
`ifndef __CAST_NETWORK_CONFIG_SVH_
`define __CAST_NETWORK_CONFIG_SVH_
`include "params.svh"
    
localparam bit [`PN-1:0] routing_table_0_0 [`PN] [`VN] = '{
'{'b00100, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_0_1 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_0_2 [`PN] [`VN] = '{
'{'b00100, 'b00000},
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_0_3 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00001, 'b00000}};

localparam bit [`PN-1:0] routing_table_0_4 [`PN] [`VN] = '{
'{'b00100, 'b00000},
'{'b00000, 'b00000},
'{'b01001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_0_5 [`PN] [`VN] = '{
'{'b10000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00001, 'b00000}};

localparam bit [`PN-1:0] routing_table_0_6 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b01001, 'b00000},
'{'b00100, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_0_7 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b10001},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_0_8 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00001},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_1_0 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00101, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_1_1 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00010, 'b00000}};

localparam bit [`PN-1:0] routing_table_1_2 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b10100, 'b00000},
'{'b01011, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_1_3 [`PN] [`VN] = '{
'{'b00100, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00001},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_1_4 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00011, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_1_5 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_1_6 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00011, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_1_7 [`PN] [`VN] = '{
'{'b00100, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00010},
'{'b00001, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_1_8 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_2_0 [`PN] [`VN] = '{
'{'b00000, 'b00100},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_2_1 [`PN] [`VN] = '{
'{'b10000, 'b00000},
'{'b00000, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_2_2 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b10101, 'b00000},
'{'b00000, 'b00000},
'{'b00010, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_2_3 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00000, 'b00011},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_2_4 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00101, 'b00000},
'{'b00010, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_2_5 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00011, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_2_6 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00011, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_2_7 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00000, 'b00010},
'{'b00001, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_2_8 [`PN] [`VN] = '{
'{'b00100, 'b00000},
'{'b00000, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_3_0 [`PN] [`VN] = '{
'{'b00100, 'b00000},
'{'b00000, 'b00101},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_3_1 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_3_2 [`PN] [`VN] = '{
'{'b00000, 'b00100},
'{'b00101, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_3_3 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00000, 'b00011},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_3_4 [`PN] [`VN] = '{
'{'b10000, 'b00000},
'{'b00101, 'b00000},
'{'b00010, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_3_5 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00011, 'b00000},
'{'b00100, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_3_6 [`PN] [`VN] = '{
'{'b01000, 'b00000},
'{'b00100, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_3_7 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00001, 'b00010},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_3_8 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_4_0 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00001},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_4_1 [`PN] [`VN] = '{
'{'b00010, 'b00000},
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_4_2 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b10001, 'b00100},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_4_3 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00001, 'b00010},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_4_4 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00101, 'b00000},
'{'b00010, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_4_5 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00011, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_4_6 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00100, 'b00000},
'{'b00011, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_4_7 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00011},
'{'b00010, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_4_8 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00010, 'b00000},
'{'b00101, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_5_0 [`PN] [`VN] = '{
'{'b00000, 'b00100},
'{'b00101, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_5_1 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_5_2 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00101},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_5_3 [`PN] [`VN] = '{
'{'b00000, 'b00010},
'{'b00100, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_5_4 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00101, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00010, 'b00000}};

localparam bit [`PN-1:0] routing_table_5_5 [`PN] [`VN] = '{
'{'b10000, 'b00000},
'{'b00100, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000},
'{'b01000, 'b00000}};

localparam bit [`PN-1:0] routing_table_5_6 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00101, 'b00000},
'{'b11000, 'b00000},
'{'b00010, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_5_7 [`PN] [`VN] = '{
'{'b10000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00010},
'{'b00101, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_5_8 [`PN] [`VN] = '{
'{'b01000, 'b00000},
'{'b00101, 'b00000},
'{'b00000, 'b00000},
'{'b00010, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_6_0 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00001, 'b00100},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_6_1 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_6_2 [`PN] [`VN] = '{
'{'b10000, 'b00000},
'{'b00000, 'b00101},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_6_3 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b10000, 'b00000},
'{'b00011, 'b00000},
'{'b00100, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_6_4 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b10000, 'b00000},
'{'b00100, 'b00000}};

localparam bit [`PN-1:0] routing_table_6_5 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b01001, 'b00000},
'{'b00010, 'b00000},
'{'b10000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_6_6 [`PN] [`VN] = '{
'{'b00000, 'b10000},
'{'b00100, 'b00000},
'{'b00000, 'b00000},
'{'b00011, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_6_7 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00101, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00010},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_6_8 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_7_0 [`PN] [`VN] = '{
'{'b10000, 'b00000},
'{'b00000, 'b00101},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_7_1 [`PN] [`VN] = '{
'{'b00010, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00101, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_7_2 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00001},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00100, 'b00000}};

localparam bit [`PN-1:0] routing_table_7_3 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b01101, 'b00000},
'{'b00010, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_7_4 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b10101, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_7_5 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00010, 'b00000},
'{'b00101, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_7_6 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00101, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_7_7 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_7_8 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_8_0 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00001},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_8_1 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_8_2 [`PN] [`VN] = '{
'{'b10000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_8_3 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00010, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_8_4 [`PN] [`VN] = '{
'{'b10000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_8_5 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000},
'{'b00010, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_8_6 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b10001, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_8_7 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00001, 'b00000},
'{'b00000, 'b00000}};

localparam bit [`PN-1:0] routing_table_8_8 [`PN] [`VN] = '{
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000},
'{'b00000, 'b00000}};

`endif
