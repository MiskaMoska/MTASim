
`ifndef                 _PARAMS_SVH_
`define                 _PARAMS_SVH_

/****************************** data width ******************************/
`define                 DW                              32

/************************** router port number **************************/
`define                 PN                              5

/************************ vc number in each port ************************/
`define                 VN                              2

/**************************** network width *****************************/
`define                 NW                              9

/**************************** network height ****************************/
`define                 NH                              9

/*************************** eject port number ***************************/
`define                 EPN                             3

`endif

