
`ifndef __CONNECTION_CONFIG_SVH_
`define __CONNECTION_CONFIG_SVH_
`include "params.svh"

localparam int cast_out_vc [`NW] [`NH] = '{
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{1, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 1, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{1, 0, 0, 1, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 1, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0}};
localparam int cast_out [`NW] [`NH] = '{
'{1, 0, 1, 0, 1, 1, 0, 0, 0},
'{0, 0, 0, 1, 0, 0, 0, 1, 0},
'{1, 1, 0, 0, 0, 0, 0, 0, 1},
'{1, 0, 1, 0, 1, 0, 1, 0, 0},
'{0, 1, 0, 0, 0, 0, 0, 0, 0},
'{1, 0, 0, 1, 0, 1, 0, 1, 1},
'{0, 0, 1, 0, 0, 0, 1, 0, 0},
'{1, 1, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 1, 0, 1, 0, 0, 0, 0}};
localparam int gather_out [`NW] [`NH] = '{
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0}};
localparam int merge_out [`NW] [`NH] = '{
'{0, 1, 0, 1, 0, 0, 1, 1, 1},
'{1, 1, 1, 0, 1, 1, 1, 0, 1},
'{0, 0, 1, 1, 1, 1, 1, 1, 0},
'{0, 1, 0, 1, 0, 1, 0, 1, 1},
'{1, 0, 1, 1, 1, 1, 1, 1, 1},
'{0, 1, 1, 0, 1, 0, 1, 0, 0},
'{1, 1, 0, 1, 1, 1, 0, 1, 1},
'{0, 0, 1, 1, 1, 1, 1, 1, 0},
'{1, 1, 0, 1, 0, 1, 1, 1, 0}};
localparam int gather_in_vc [`NW] [`NH] = '{
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0}};
localparam int merge_in [`NW] [`NH] = '{
'{0, 0, 1, 0, 1, 0, 0, 0, 0},
'{0, 0, 0, 1, 0, 0, 0, 1, 0},
'{1, 1, 0, 0, 0, 0, 0, 0, 1},
'{1, 0, 1, 0, 1, 0, 1, 0, 0},
'{0, 1, 0, 0, 0, 0, 0, 0, 0},
'{1, 0, 0, 1, 0, 1, 0, 1, 1},
'{0, 0, 1, 0, 0, 0, 1, 0, 0},
'{1, 1, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 1, 0, 1, 0, 0, 0, 0}};
localparam int gather_out_vc [`NW] [`NH] = '{
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0}};
localparam int cast_in_vc [`NW] [`NH] = '{
'{0, 0, 0, 0, 0, 0, 0, 1, 1},
'{0, 0, 0, 1, 0, 0, 0, 0, 0},
'{0, 0, 0, 1, 0, 0, 0, 0, 0},
'{1, 0, 0, 1, 0, 0, 0, 0, 0},
'{1, 0, 0, 0, 0, 0, 0, 1, 0},
'{0, 0, 1, 0, 0, 0, 0, 0, 0},
'{0, 0, 1, 0, 0, 0, 0, 0, 0},
'{1, 0, 1, 0, 0, 0, 0, 0, 0},
'{1, 0, 0, 0, 0, 0, 0, 0, 0}};
localparam int gather_in [`NW] [`NH] = '{
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0},
'{0, 0, 0, 0, 0, 0, 0, 0, 0}};

`endif

