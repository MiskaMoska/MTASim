`ifndef     __PARAMS_SVH__
`define     __PARAMS_SVH__

`define     QW          32
`define     XH          1152
`define     XW          256

`endif