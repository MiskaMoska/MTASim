
//Cast Network
//Width: 6
//Height:8

`include "params.svh"
`include "cast_network_config.svh"

module cast_network(
    input       wire                            clk,
    input       wire                            rstn,

    input       wire        [`VN-1:0]           vc_i [`NW] [`NH],
    input       wire        [`DW-1:0]           data_i [`NW] [`NH],
    input       wire                            valid_i [`NW] [`NH],
    output      reg                             ready_o [`NW] [`NH],

    output      reg         [`VN-1:0]           vc_o [`NW] [`NH],
    output      reg         [`DW-1:0]           data_o [`NW] [`NH],
    output      reg                             valid_o [`NW] [`NH],
    input       wire                            ready_i [`NW] [`NH]
);

logic [`VN-1:0] vc_i_0_0[5];
logic [`DW-1:0] data_i_0_0[5];
logic valid_i_0_0[5], ready_i_0_0[5];    
logic [`VN-1:0] vc_o_0_0[5];
logic [`DW-1:0] data_o_0_0[5];
logic valid_o_0_0[5], ready_o_0_0[5];        

logic [`VN-1:0] vc_i_0_1[5];
logic [`DW-1:0] data_i_0_1[5];
logic valid_i_0_1[5], ready_i_0_1[5];    
logic [`VN-1:0] vc_o_0_1[5];
logic [`DW-1:0] data_o_0_1[5];
logic valid_o_0_1[5], ready_o_0_1[5];        

logic [`VN-1:0] vc_i_0_2[5];
logic [`DW-1:0] data_i_0_2[5];
logic valid_i_0_2[5], ready_i_0_2[5];    
logic [`VN-1:0] vc_o_0_2[5];
logic [`DW-1:0] data_o_0_2[5];
logic valid_o_0_2[5], ready_o_0_2[5];        

logic [`VN-1:0] vc_i_0_3[5];
logic [`DW-1:0] data_i_0_3[5];
logic valid_i_0_3[5], ready_i_0_3[5];    
logic [`VN-1:0] vc_o_0_3[5];
logic [`DW-1:0] data_o_0_3[5];
logic valid_o_0_3[5], ready_o_0_3[5];        

logic [`VN-1:0] vc_i_0_4[5];
logic [`DW-1:0] data_i_0_4[5];
logic valid_i_0_4[5], ready_i_0_4[5];    
logic [`VN-1:0] vc_o_0_4[5];
logic [`DW-1:0] data_o_0_4[5];
logic valid_o_0_4[5], ready_o_0_4[5];        

logic [`VN-1:0] vc_i_0_5[5];
logic [`DW-1:0] data_i_0_5[5];
logic valid_i_0_5[5], ready_i_0_5[5];    
logic [`VN-1:0] vc_o_0_5[5];
logic [`DW-1:0] data_o_0_5[5];
logic valid_o_0_5[5], ready_o_0_5[5];        

logic [`VN-1:0] vc_i_0_6[5];
logic [`DW-1:0] data_i_0_6[5];
logic valid_i_0_6[5], ready_i_0_6[5];    
logic [`VN-1:0] vc_o_0_6[5];
logic [`DW-1:0] data_o_0_6[5];
logic valid_o_0_6[5], ready_o_0_6[5];        

logic [`VN-1:0] vc_i_0_7[5];
logic [`DW-1:0] data_i_0_7[5];
logic valid_i_0_7[5], ready_i_0_7[5];    
logic [`VN-1:0] vc_o_0_7[5];
logic [`DW-1:0] data_o_0_7[5];
logic valid_o_0_7[5], ready_o_0_7[5];        

logic [`VN-1:0] vc_i_1_0[5];
logic [`DW-1:0] data_i_1_0[5];
logic valid_i_1_0[5], ready_i_1_0[5];    
logic [`VN-1:0] vc_o_1_0[5];
logic [`DW-1:0] data_o_1_0[5];
logic valid_o_1_0[5], ready_o_1_0[5];        

logic [`VN-1:0] vc_i_1_1[5];
logic [`DW-1:0] data_i_1_1[5];
logic valid_i_1_1[5], ready_i_1_1[5];    
logic [`VN-1:0] vc_o_1_1[5];
logic [`DW-1:0] data_o_1_1[5];
logic valid_o_1_1[5], ready_o_1_1[5];        

logic [`VN-1:0] vc_i_1_2[5];
logic [`DW-1:0] data_i_1_2[5];
logic valid_i_1_2[5], ready_i_1_2[5];    
logic [`VN-1:0] vc_o_1_2[5];
logic [`DW-1:0] data_o_1_2[5];
logic valid_o_1_2[5], ready_o_1_2[5];        

logic [`VN-1:0] vc_i_1_3[5];
logic [`DW-1:0] data_i_1_3[5];
logic valid_i_1_3[5], ready_i_1_3[5];    
logic [`VN-1:0] vc_o_1_3[5];
logic [`DW-1:0] data_o_1_3[5];
logic valid_o_1_3[5], ready_o_1_3[5];        

logic [`VN-1:0] vc_i_1_4[5];
logic [`DW-1:0] data_i_1_4[5];
logic valid_i_1_4[5], ready_i_1_4[5];    
logic [`VN-1:0] vc_o_1_4[5];
logic [`DW-1:0] data_o_1_4[5];
logic valid_o_1_4[5], ready_o_1_4[5];        

logic [`VN-1:0] vc_i_1_5[5];
logic [`DW-1:0] data_i_1_5[5];
logic valid_i_1_5[5], ready_i_1_5[5];    
logic [`VN-1:0] vc_o_1_5[5];
logic [`DW-1:0] data_o_1_5[5];
logic valid_o_1_5[5], ready_o_1_5[5];        

logic [`VN-1:0] vc_i_1_6[5];
logic [`DW-1:0] data_i_1_6[5];
logic valid_i_1_6[5], ready_i_1_6[5];    
logic [`VN-1:0] vc_o_1_6[5];
logic [`DW-1:0] data_o_1_6[5];
logic valid_o_1_6[5], ready_o_1_6[5];        

logic [`VN-1:0] vc_i_1_7[5];
logic [`DW-1:0] data_i_1_7[5];
logic valid_i_1_7[5], ready_i_1_7[5];    
logic [`VN-1:0] vc_o_1_7[5];
logic [`DW-1:0] data_o_1_7[5];
logic valid_o_1_7[5], ready_o_1_7[5];        

logic [`VN-1:0] vc_i_2_0[5];
logic [`DW-1:0] data_i_2_0[5];
logic valid_i_2_0[5], ready_i_2_0[5];    
logic [`VN-1:0] vc_o_2_0[5];
logic [`DW-1:0] data_o_2_0[5];
logic valid_o_2_0[5], ready_o_2_0[5];        

logic [`VN-1:0] vc_i_2_1[5];
logic [`DW-1:0] data_i_2_1[5];
logic valid_i_2_1[5], ready_i_2_1[5];    
logic [`VN-1:0] vc_o_2_1[5];
logic [`DW-1:0] data_o_2_1[5];
logic valid_o_2_1[5], ready_o_2_1[5];        

logic [`VN-1:0] vc_i_2_2[5];
logic [`DW-1:0] data_i_2_2[5];
logic valid_i_2_2[5], ready_i_2_2[5];    
logic [`VN-1:0] vc_o_2_2[5];
logic [`DW-1:0] data_o_2_2[5];
logic valid_o_2_2[5], ready_o_2_2[5];        

logic [`VN-1:0] vc_i_2_3[5];
logic [`DW-1:0] data_i_2_3[5];
logic valid_i_2_3[5], ready_i_2_3[5];    
logic [`VN-1:0] vc_o_2_3[5];
logic [`DW-1:0] data_o_2_3[5];
logic valid_o_2_3[5], ready_o_2_3[5];        

logic [`VN-1:0] vc_i_2_4[5];
logic [`DW-1:0] data_i_2_4[5];
logic valid_i_2_4[5], ready_i_2_4[5];    
logic [`VN-1:0] vc_o_2_4[5];
logic [`DW-1:0] data_o_2_4[5];
logic valid_o_2_4[5], ready_o_2_4[5];        

logic [`VN-1:0] vc_i_2_5[5];
logic [`DW-1:0] data_i_2_5[5];
logic valid_i_2_5[5], ready_i_2_5[5];    
logic [`VN-1:0] vc_o_2_5[5];
logic [`DW-1:0] data_o_2_5[5];
logic valid_o_2_5[5], ready_o_2_5[5];        

logic [`VN-1:0] vc_i_2_6[5];
logic [`DW-1:0] data_i_2_6[5];
logic valid_i_2_6[5], ready_i_2_6[5];    
logic [`VN-1:0] vc_o_2_6[5];
logic [`DW-1:0] data_o_2_6[5];
logic valid_o_2_6[5], ready_o_2_6[5];        

logic [`VN-1:0] vc_i_2_7[5];
logic [`DW-1:0] data_i_2_7[5];
logic valid_i_2_7[5], ready_i_2_7[5];    
logic [`VN-1:0] vc_o_2_7[5];
logic [`DW-1:0] data_o_2_7[5];
logic valid_o_2_7[5], ready_o_2_7[5];        

logic [`VN-1:0] vc_i_3_0[5];
logic [`DW-1:0] data_i_3_0[5];
logic valid_i_3_0[5], ready_i_3_0[5];    
logic [`VN-1:0] vc_o_3_0[5];
logic [`DW-1:0] data_o_3_0[5];
logic valid_o_3_0[5], ready_o_3_0[5];        

logic [`VN-1:0] vc_i_3_1[5];
logic [`DW-1:0] data_i_3_1[5];
logic valid_i_3_1[5], ready_i_3_1[5];    
logic [`VN-1:0] vc_o_3_1[5];
logic [`DW-1:0] data_o_3_1[5];
logic valid_o_3_1[5], ready_o_3_1[5];        

logic [`VN-1:0] vc_i_3_2[5];
logic [`DW-1:0] data_i_3_2[5];
logic valid_i_3_2[5], ready_i_3_2[5];    
logic [`VN-1:0] vc_o_3_2[5];
logic [`DW-1:0] data_o_3_2[5];
logic valid_o_3_2[5], ready_o_3_2[5];        

logic [`VN-1:0] vc_i_3_3[5];
logic [`DW-1:0] data_i_3_3[5];
logic valid_i_3_3[5], ready_i_3_3[5];    
logic [`VN-1:0] vc_o_3_3[5];
logic [`DW-1:0] data_o_3_3[5];
logic valid_o_3_3[5], ready_o_3_3[5];        

logic [`VN-1:0] vc_i_3_4[5];
logic [`DW-1:0] data_i_3_4[5];
logic valid_i_3_4[5], ready_i_3_4[5];    
logic [`VN-1:0] vc_o_3_4[5];
logic [`DW-1:0] data_o_3_4[5];
logic valid_o_3_4[5], ready_o_3_4[5];        

logic [`VN-1:0] vc_i_3_5[5];
logic [`DW-1:0] data_i_3_5[5];
logic valid_i_3_5[5], ready_i_3_5[5];    
logic [`VN-1:0] vc_o_3_5[5];
logic [`DW-1:0] data_o_3_5[5];
logic valid_o_3_5[5], ready_o_3_5[5];        

logic [`VN-1:0] vc_i_3_6[5];
logic [`DW-1:0] data_i_3_6[5];
logic valid_i_3_6[5], ready_i_3_6[5];    
logic [`VN-1:0] vc_o_3_6[5];
logic [`DW-1:0] data_o_3_6[5];
logic valid_o_3_6[5], ready_o_3_6[5];        

logic [`VN-1:0] vc_i_3_7[5];
logic [`DW-1:0] data_i_3_7[5];
logic valid_i_3_7[5], ready_i_3_7[5];    
logic [`VN-1:0] vc_o_3_7[5];
logic [`DW-1:0] data_o_3_7[5];
logic valid_o_3_7[5], ready_o_3_7[5];        

logic [`VN-1:0] vc_i_4_0[5];
logic [`DW-1:0] data_i_4_0[5];
logic valid_i_4_0[5], ready_i_4_0[5];    
logic [`VN-1:0] vc_o_4_0[5];
logic [`DW-1:0] data_o_4_0[5];
logic valid_o_4_0[5], ready_o_4_0[5];        

logic [`VN-1:0] vc_i_4_1[5];
logic [`DW-1:0] data_i_4_1[5];
logic valid_i_4_1[5], ready_i_4_1[5];    
logic [`VN-1:0] vc_o_4_1[5];
logic [`DW-1:0] data_o_4_1[5];
logic valid_o_4_1[5], ready_o_4_1[5];        

logic [`VN-1:0] vc_i_4_2[5];
logic [`DW-1:0] data_i_4_2[5];
logic valid_i_4_2[5], ready_i_4_2[5];    
logic [`VN-1:0] vc_o_4_2[5];
logic [`DW-1:0] data_o_4_2[5];
logic valid_o_4_2[5], ready_o_4_2[5];        

logic [`VN-1:0] vc_i_4_3[5];
logic [`DW-1:0] data_i_4_3[5];
logic valid_i_4_3[5], ready_i_4_3[5];    
logic [`VN-1:0] vc_o_4_3[5];
logic [`DW-1:0] data_o_4_3[5];
logic valid_o_4_3[5], ready_o_4_3[5];        

logic [`VN-1:0] vc_i_4_4[5];
logic [`DW-1:0] data_i_4_4[5];
logic valid_i_4_4[5], ready_i_4_4[5];    
logic [`VN-1:0] vc_o_4_4[5];
logic [`DW-1:0] data_o_4_4[5];
logic valid_o_4_4[5], ready_o_4_4[5];        

logic [`VN-1:0] vc_i_4_5[5];
logic [`DW-1:0] data_i_4_5[5];
logic valid_i_4_5[5], ready_i_4_5[5];    
logic [`VN-1:0] vc_o_4_5[5];
logic [`DW-1:0] data_o_4_5[5];
logic valid_o_4_5[5], ready_o_4_5[5];        

logic [`VN-1:0] vc_i_4_6[5];
logic [`DW-1:0] data_i_4_6[5];
logic valid_i_4_6[5], ready_i_4_6[5];    
logic [`VN-1:0] vc_o_4_6[5];
logic [`DW-1:0] data_o_4_6[5];
logic valid_o_4_6[5], ready_o_4_6[5];        

logic [`VN-1:0] vc_i_4_7[5];
logic [`DW-1:0] data_i_4_7[5];
logic valid_i_4_7[5], ready_i_4_7[5];    
logic [`VN-1:0] vc_o_4_7[5];
logic [`DW-1:0] data_o_4_7[5];
logic valid_o_4_7[5], ready_o_4_7[5];        

logic [`VN-1:0] vc_i_5_0[5];
logic [`DW-1:0] data_i_5_0[5];
logic valid_i_5_0[5], ready_i_5_0[5];    
logic [`VN-1:0] vc_o_5_0[5];
logic [`DW-1:0] data_o_5_0[5];
logic valid_o_5_0[5], ready_o_5_0[5];        

logic [`VN-1:0] vc_i_5_1[5];
logic [`DW-1:0] data_i_5_1[5];
logic valid_i_5_1[5], ready_i_5_1[5];    
logic [`VN-1:0] vc_o_5_1[5];
logic [`DW-1:0] data_o_5_1[5];
logic valid_o_5_1[5], ready_o_5_1[5];        

logic [`VN-1:0] vc_i_5_2[5];
logic [`DW-1:0] data_i_5_2[5];
logic valid_i_5_2[5], ready_i_5_2[5];    
logic [`VN-1:0] vc_o_5_2[5];
logic [`DW-1:0] data_o_5_2[5];
logic valid_o_5_2[5], ready_o_5_2[5];        

logic [`VN-1:0] vc_i_5_3[5];
logic [`DW-1:0] data_i_5_3[5];
logic valid_i_5_3[5], ready_i_5_3[5];    
logic [`VN-1:0] vc_o_5_3[5];
logic [`DW-1:0] data_o_5_3[5];
logic valid_o_5_3[5], ready_o_5_3[5];        

logic [`VN-1:0] vc_i_5_4[5];
logic [`DW-1:0] data_i_5_4[5];
logic valid_i_5_4[5], ready_i_5_4[5];    
logic [`VN-1:0] vc_o_5_4[5];
logic [`DW-1:0] data_o_5_4[5];
logic valid_o_5_4[5], ready_o_5_4[5];        

logic [`VN-1:0] vc_i_5_5[5];
logic [`DW-1:0] data_i_5_5[5];
logic valid_i_5_5[5], ready_i_5_5[5];    
logic [`VN-1:0] vc_o_5_5[5];
logic [`DW-1:0] data_o_5_5[5];
logic valid_o_5_5[5], ready_o_5_5[5];        

logic [`VN-1:0] vc_i_5_6[5];
logic [`DW-1:0] data_i_5_6[5];
logic valid_i_5_6[5], ready_i_5_6[5];    
logic [`VN-1:0] vc_o_5_6[5];
logic [`DW-1:0] data_o_5_6[5];
logic valid_o_5_6[5], ready_o_5_6[5];        

logic [`VN-1:0] vc_i_5_7[5];
logic [`DW-1:0] data_i_5_7[5];
logic valid_i_5_7[5], ready_i_5_7[5];    
logic [`VN-1:0] vc_o_5_7[5];
logic [`DW-1:0] data_o_5_7[5];
logic valid_o_5_7[5], ready_o_5_7[5];        

always_comb begin
    vc_o[0][0] = vc_o_0_0[0];
    data_o[0][0] = data_o_0_0[0];
    valid_o[0][0] = valid_o_0_0[0];
    ready_o[0][0] = ready_o_0_0[0];
    vc_o[0][1] = vc_o_0_1[0];
    data_o[0][1] = data_o_0_1[0];
    valid_o[0][1] = valid_o_0_1[0];
    ready_o[0][1] = ready_o_0_1[0];
    vc_o[0][2] = vc_o_0_2[0];
    data_o[0][2] = data_o_0_2[0];
    valid_o[0][2] = valid_o_0_2[0];
    ready_o[0][2] = ready_o_0_2[0];
    vc_o[0][3] = vc_o_0_3[0];
    data_o[0][3] = data_o_0_3[0];
    valid_o[0][3] = valid_o_0_3[0];
    ready_o[0][3] = ready_o_0_3[0];
    vc_o[0][4] = vc_o_0_4[0];
    data_o[0][4] = data_o_0_4[0];
    valid_o[0][4] = valid_o_0_4[0];
    ready_o[0][4] = ready_o_0_4[0];
    vc_o[0][5] = vc_o_0_5[0];
    data_o[0][5] = data_o_0_5[0];
    valid_o[0][5] = valid_o_0_5[0];
    ready_o[0][5] = ready_o_0_5[0];
    vc_o[0][6] = vc_o_0_6[0];
    data_o[0][6] = data_o_0_6[0];
    valid_o[0][6] = valid_o_0_6[0];
    ready_o[0][6] = ready_o_0_6[0];
    vc_o[0][7] = vc_o_0_7[0];
    data_o[0][7] = data_o_0_7[0];
    valid_o[0][7] = valid_o_0_7[0];
    ready_o[0][7] = ready_o_0_7[0];
    vc_o[1][0] = vc_o_1_0[0];
    data_o[1][0] = data_o_1_0[0];
    valid_o[1][0] = valid_o_1_0[0];
    ready_o[1][0] = ready_o_1_0[0];
    vc_o[1][1] = vc_o_1_1[0];
    data_o[1][1] = data_o_1_1[0];
    valid_o[1][1] = valid_o_1_1[0];
    ready_o[1][1] = ready_o_1_1[0];
    vc_o[1][2] = vc_o_1_2[0];
    data_o[1][2] = data_o_1_2[0];
    valid_o[1][2] = valid_o_1_2[0];
    ready_o[1][2] = ready_o_1_2[0];
    vc_o[1][3] = vc_o_1_3[0];
    data_o[1][3] = data_o_1_3[0];
    valid_o[1][3] = valid_o_1_3[0];
    ready_o[1][3] = ready_o_1_3[0];
    vc_o[1][4] = vc_o_1_4[0];
    data_o[1][4] = data_o_1_4[0];
    valid_o[1][4] = valid_o_1_4[0];
    ready_o[1][4] = ready_o_1_4[0];
    vc_o[1][5] = vc_o_1_5[0];
    data_o[1][5] = data_o_1_5[0];
    valid_o[1][5] = valid_o_1_5[0];
    ready_o[1][5] = ready_o_1_5[0];
    vc_o[1][6] = vc_o_1_6[0];
    data_o[1][6] = data_o_1_6[0];
    valid_o[1][6] = valid_o_1_6[0];
    ready_o[1][6] = ready_o_1_6[0];
    vc_o[1][7] = vc_o_1_7[0];
    data_o[1][7] = data_o_1_7[0];
    valid_o[1][7] = valid_o_1_7[0];
    ready_o[1][7] = ready_o_1_7[0];
    vc_o[2][0] = vc_o_2_0[0];
    data_o[2][0] = data_o_2_0[0];
    valid_o[2][0] = valid_o_2_0[0];
    ready_o[2][0] = ready_o_2_0[0];
    vc_o[2][1] = vc_o_2_1[0];
    data_o[2][1] = data_o_2_1[0];
    valid_o[2][1] = valid_o_2_1[0];
    ready_o[2][1] = ready_o_2_1[0];
    vc_o[2][2] = vc_o_2_2[0];
    data_o[2][2] = data_o_2_2[0];
    valid_o[2][2] = valid_o_2_2[0];
    ready_o[2][2] = ready_o_2_2[0];
    vc_o[2][3] = vc_o_2_3[0];
    data_o[2][3] = data_o_2_3[0];
    valid_o[2][3] = valid_o_2_3[0];
    ready_o[2][3] = ready_o_2_3[0];
    vc_o[2][4] = vc_o_2_4[0];
    data_o[2][4] = data_o_2_4[0];
    valid_o[2][4] = valid_o_2_4[0];
    ready_o[2][4] = ready_o_2_4[0];
    vc_o[2][5] = vc_o_2_5[0];
    data_o[2][5] = data_o_2_5[0];
    valid_o[2][5] = valid_o_2_5[0];
    ready_o[2][5] = ready_o_2_5[0];
    vc_o[2][6] = vc_o_2_6[0];
    data_o[2][6] = data_o_2_6[0];
    valid_o[2][6] = valid_o_2_6[0];
    ready_o[2][6] = ready_o_2_6[0];
    vc_o[2][7] = vc_o_2_7[0];
    data_o[2][7] = data_o_2_7[0];
    valid_o[2][7] = valid_o_2_7[0];
    ready_o[2][7] = ready_o_2_7[0];
    vc_o[3][0] = vc_o_3_0[0];
    data_o[3][0] = data_o_3_0[0];
    valid_o[3][0] = valid_o_3_0[0];
    ready_o[3][0] = ready_o_3_0[0];
    vc_o[3][1] = vc_o_3_1[0];
    data_o[3][1] = data_o_3_1[0];
    valid_o[3][1] = valid_o_3_1[0];
    ready_o[3][1] = ready_o_3_1[0];
    vc_o[3][2] = vc_o_3_2[0];
    data_o[3][2] = data_o_3_2[0];
    valid_o[3][2] = valid_o_3_2[0];
    ready_o[3][2] = ready_o_3_2[0];
    vc_o[3][3] = vc_o_3_3[0];
    data_o[3][3] = data_o_3_3[0];
    valid_o[3][3] = valid_o_3_3[0];
    ready_o[3][3] = ready_o_3_3[0];
    vc_o[3][4] = vc_o_3_4[0];
    data_o[3][4] = data_o_3_4[0];
    valid_o[3][4] = valid_o_3_4[0];
    ready_o[3][4] = ready_o_3_4[0];
    vc_o[3][5] = vc_o_3_5[0];
    data_o[3][5] = data_o_3_5[0];
    valid_o[3][5] = valid_o_3_5[0];
    ready_o[3][5] = ready_o_3_5[0];
    vc_o[3][6] = vc_o_3_6[0];
    data_o[3][6] = data_o_3_6[0];
    valid_o[3][6] = valid_o_3_6[0];
    ready_o[3][6] = ready_o_3_6[0];
    vc_o[3][7] = vc_o_3_7[0];
    data_o[3][7] = data_o_3_7[0];
    valid_o[3][7] = valid_o_3_7[0];
    ready_o[3][7] = ready_o_3_7[0];
    vc_o[4][0] = vc_o_4_0[0];
    data_o[4][0] = data_o_4_0[0];
    valid_o[4][0] = valid_o_4_0[0];
    ready_o[4][0] = ready_o_4_0[0];
    vc_o[4][1] = vc_o_4_1[0];
    data_o[4][1] = data_o_4_1[0];
    valid_o[4][1] = valid_o_4_1[0];
    ready_o[4][1] = ready_o_4_1[0];
    vc_o[4][2] = vc_o_4_2[0];
    data_o[4][2] = data_o_4_2[0];
    valid_o[4][2] = valid_o_4_2[0];
    ready_o[4][2] = ready_o_4_2[0];
    vc_o[4][3] = vc_o_4_3[0];
    data_o[4][3] = data_o_4_3[0];
    valid_o[4][3] = valid_o_4_3[0];
    ready_o[4][3] = ready_o_4_3[0];
    vc_o[4][4] = vc_o_4_4[0];
    data_o[4][4] = data_o_4_4[0];
    valid_o[4][4] = valid_o_4_4[0];
    ready_o[4][4] = ready_o_4_4[0];
    vc_o[4][5] = vc_o_4_5[0];
    data_o[4][5] = data_o_4_5[0];
    valid_o[4][5] = valid_o_4_5[0];
    ready_o[4][5] = ready_o_4_5[0];
    vc_o[4][6] = vc_o_4_6[0];
    data_o[4][6] = data_o_4_6[0];
    valid_o[4][6] = valid_o_4_6[0];
    ready_o[4][6] = ready_o_4_6[0];
    vc_o[4][7] = vc_o_4_7[0];
    data_o[4][7] = data_o_4_7[0];
    valid_o[4][7] = valid_o_4_7[0];
    ready_o[4][7] = ready_o_4_7[0];
    vc_o[5][0] = vc_o_5_0[0];
    data_o[5][0] = data_o_5_0[0];
    valid_o[5][0] = valid_o_5_0[0];
    ready_o[5][0] = ready_o_5_0[0];
    vc_o[5][1] = vc_o_5_1[0];
    data_o[5][1] = data_o_5_1[0];
    valid_o[5][1] = valid_o_5_1[0];
    ready_o[5][1] = ready_o_5_1[0];
    vc_o[5][2] = vc_o_5_2[0];
    data_o[5][2] = data_o_5_2[0];
    valid_o[5][2] = valid_o_5_2[0];
    ready_o[5][2] = ready_o_5_2[0];
    vc_o[5][3] = vc_o_5_3[0];
    data_o[5][3] = data_o_5_3[0];
    valid_o[5][3] = valid_o_5_3[0];
    ready_o[5][3] = ready_o_5_3[0];
    vc_o[5][4] = vc_o_5_4[0];
    data_o[5][4] = data_o_5_4[0];
    valid_o[5][4] = valid_o_5_4[0];
    ready_o[5][4] = ready_o_5_4[0];
    vc_o[5][5] = vc_o_5_5[0];
    data_o[5][5] = data_o_5_5[0];
    valid_o[5][5] = valid_o_5_5[0];
    ready_o[5][5] = ready_o_5_5[0];
    vc_o[5][6] = vc_o_5_6[0];
    data_o[5][6] = data_o_5_6[0];
    valid_o[5][6] = valid_o_5_6[0];
    ready_o[5][6] = ready_o_5_6[0];
    vc_o[5][7] = vc_o_5_7[0];
    data_o[5][7] = data_o_5_7[0];
    valid_o[5][7] = valid_o_5_7[0];
    ready_o[5][7] = ready_o_5_7[0];
end

/*Router 0,0*/    
cast_router #(
    .routing_table                  (routing_table_0_0)
)router_0_0(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_0_0),
    .data_i                         (data_i_0_0),
    .valid_i                        (valid_i_0_0),
    .ready_o                        (ready_o_0_0),
    .vc_o                           (vc_o_0_0),
    .data_o                         (data_o_0_0),
    .valid_o                        (valid_o_0_0),
    .ready_i                        (ready_i_0_0)
);


always_comb begin
    vc_i_0_0[4] = vc_o_0_1[3];
    data_i_0_0[4] = data_o_0_1[3];
    valid_i_0_0[4] = valid_o_0_1[3];
    ready_i_0_0[4] = ready_o_0_1[3];
    vc_i_0_0[2] = vc_o_1_0[1];
    data_i_0_0[2] = data_o_1_0[1];
    valid_i_0_0[2] = valid_o_1_0[1];
    ready_i_0_0[2] = ready_o_1_0[1];
    vc_i_0_0[0] = vc_i[0][0];
    data_i_0_0[0] = data_i[0][0];
    valid_i_0_0[0] = valid_i[0][0];
    ready_i_0_0[0] = ready_i[0][0];
end


/*Router 0,1*/    
cast_router #(
    .routing_table                  (routing_table_0_1)
)router_0_1(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_0_1),
    .data_i                         (data_i_0_1),
    .valid_i                        (valid_i_0_1),
    .ready_o                        (ready_o_0_1),
    .vc_o                           (vc_o_0_1),
    .data_o                         (data_o_0_1),
    .valid_o                        (valid_o_0_1),
    .ready_i                        (ready_i_0_1)
);


always_comb begin
    vc_i_0_1[3] = vc_o_0_0[4];
    data_i_0_1[3] = data_o_0_0[4];
    valid_i_0_1[3] = valid_o_0_0[4];
    ready_i_0_1[3] = ready_o_0_0[4];
    vc_i_0_1[4] = vc_o_0_2[3];
    data_i_0_1[4] = data_o_0_2[3];
    valid_i_0_1[4] = valid_o_0_2[3];
    ready_i_0_1[4] = ready_o_0_2[3];
    vc_i_0_1[2] = vc_o_1_1[1];
    data_i_0_1[2] = data_o_1_1[1];
    valid_i_0_1[2] = valid_o_1_1[1];
    ready_i_0_1[2] = ready_o_1_1[1];
    vc_i_0_1[0] = vc_i[0][1];
    data_i_0_1[0] = data_i[0][1];
    valid_i_0_1[0] = valid_i[0][1];
    ready_i_0_1[0] = ready_i[0][1];
end


/*Router 0,2*/    
cast_router #(
    .routing_table                  (routing_table_0_2)
)router_0_2(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_0_2),
    .data_i                         (data_i_0_2),
    .valid_i                        (valid_i_0_2),
    .ready_o                        (ready_o_0_2),
    .vc_o                           (vc_o_0_2),
    .data_o                         (data_o_0_2),
    .valid_o                        (valid_o_0_2),
    .ready_i                        (ready_i_0_2)
);


always_comb begin
    vc_i_0_2[3] = vc_o_0_1[4];
    data_i_0_2[3] = data_o_0_1[4];
    valid_i_0_2[3] = valid_o_0_1[4];
    ready_i_0_2[3] = ready_o_0_1[4];
    vc_i_0_2[4] = vc_o_0_3[3];
    data_i_0_2[4] = data_o_0_3[3];
    valid_i_0_2[4] = valid_o_0_3[3];
    ready_i_0_2[4] = ready_o_0_3[3];
    vc_i_0_2[2] = vc_o_1_2[1];
    data_i_0_2[2] = data_o_1_2[1];
    valid_i_0_2[2] = valid_o_1_2[1];
    ready_i_0_2[2] = ready_o_1_2[1];
    vc_i_0_2[0] = vc_i[0][2];
    data_i_0_2[0] = data_i[0][2];
    valid_i_0_2[0] = valid_i[0][2];
    ready_i_0_2[0] = ready_i[0][2];
end


/*Router 0,3*/    
cast_router #(
    .routing_table                  (routing_table_0_3)
)router_0_3(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_0_3),
    .data_i                         (data_i_0_3),
    .valid_i                        (valid_i_0_3),
    .ready_o                        (ready_o_0_3),
    .vc_o                           (vc_o_0_3),
    .data_o                         (data_o_0_3),
    .valid_o                        (valid_o_0_3),
    .ready_i                        (ready_i_0_3)
);


always_comb begin
    vc_i_0_3[3] = vc_o_0_2[4];
    data_i_0_3[3] = data_o_0_2[4];
    valid_i_0_3[3] = valid_o_0_2[4];
    ready_i_0_3[3] = ready_o_0_2[4];
    vc_i_0_3[4] = vc_o_0_4[3];
    data_i_0_3[4] = data_o_0_4[3];
    valid_i_0_3[4] = valid_o_0_4[3];
    ready_i_0_3[4] = ready_o_0_4[3];
    vc_i_0_3[2] = vc_o_1_3[1];
    data_i_0_3[2] = data_o_1_3[1];
    valid_i_0_3[2] = valid_o_1_3[1];
    ready_i_0_3[2] = ready_o_1_3[1];
    vc_i_0_3[0] = vc_i[0][3];
    data_i_0_3[0] = data_i[0][3];
    valid_i_0_3[0] = valid_i[0][3];
    ready_i_0_3[0] = ready_i[0][3];
end


/*Router 0,4*/    
cast_router #(
    .routing_table                  (routing_table_0_4)
)router_0_4(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_0_4),
    .data_i                         (data_i_0_4),
    .valid_i                        (valid_i_0_4),
    .ready_o                        (ready_o_0_4),
    .vc_o                           (vc_o_0_4),
    .data_o                         (data_o_0_4),
    .valid_o                        (valid_o_0_4),
    .ready_i                        (ready_i_0_4)
);


always_comb begin
    vc_i_0_4[3] = vc_o_0_3[4];
    data_i_0_4[3] = data_o_0_3[4];
    valid_i_0_4[3] = valid_o_0_3[4];
    ready_i_0_4[3] = ready_o_0_3[4];
    vc_i_0_4[4] = vc_o_0_5[3];
    data_i_0_4[4] = data_o_0_5[3];
    valid_i_0_4[4] = valid_o_0_5[3];
    ready_i_0_4[4] = ready_o_0_5[3];
    vc_i_0_4[2] = vc_o_1_4[1];
    data_i_0_4[2] = data_o_1_4[1];
    valid_i_0_4[2] = valid_o_1_4[1];
    ready_i_0_4[2] = ready_o_1_4[1];
    vc_i_0_4[0] = vc_i[0][4];
    data_i_0_4[0] = data_i[0][4];
    valid_i_0_4[0] = valid_i[0][4];
    ready_i_0_4[0] = ready_i[0][4];
end


/*Router 0,5*/    
cast_router #(
    .routing_table                  (routing_table_0_5)
)router_0_5(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_0_5),
    .data_i                         (data_i_0_5),
    .valid_i                        (valid_i_0_5),
    .ready_o                        (ready_o_0_5),
    .vc_o                           (vc_o_0_5),
    .data_o                         (data_o_0_5),
    .valid_o                        (valid_o_0_5),
    .ready_i                        (ready_i_0_5)
);


always_comb begin
    vc_i_0_5[3] = vc_o_0_4[4];
    data_i_0_5[3] = data_o_0_4[4];
    valid_i_0_5[3] = valid_o_0_4[4];
    ready_i_0_5[3] = ready_o_0_4[4];
    vc_i_0_5[4] = vc_o_0_6[3];
    data_i_0_5[4] = data_o_0_6[3];
    valid_i_0_5[4] = valid_o_0_6[3];
    ready_i_0_5[4] = ready_o_0_6[3];
    vc_i_0_5[2] = vc_o_1_5[1];
    data_i_0_5[2] = data_o_1_5[1];
    valid_i_0_5[2] = valid_o_1_5[1];
    ready_i_0_5[2] = ready_o_1_5[1];
    vc_i_0_5[0] = vc_i[0][5];
    data_i_0_5[0] = data_i[0][5];
    valid_i_0_5[0] = valid_i[0][5];
    ready_i_0_5[0] = ready_i[0][5];
end


/*Router 0,6*/    
cast_router #(
    .routing_table                  (routing_table_0_6)
)router_0_6(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_0_6),
    .data_i                         (data_i_0_6),
    .valid_i                        (valid_i_0_6),
    .ready_o                        (ready_o_0_6),
    .vc_o                           (vc_o_0_6),
    .data_o                         (data_o_0_6),
    .valid_o                        (valid_o_0_6),
    .ready_i                        (ready_i_0_6)
);


always_comb begin
    vc_i_0_6[3] = vc_o_0_5[4];
    data_i_0_6[3] = data_o_0_5[4];
    valid_i_0_6[3] = valid_o_0_5[4];
    ready_i_0_6[3] = ready_o_0_5[4];
    vc_i_0_6[4] = vc_o_0_7[3];
    data_i_0_6[4] = data_o_0_7[3];
    valid_i_0_6[4] = valid_o_0_7[3];
    ready_i_0_6[4] = ready_o_0_7[3];
    vc_i_0_6[2] = vc_o_1_6[1];
    data_i_0_6[2] = data_o_1_6[1];
    valid_i_0_6[2] = valid_o_1_6[1];
    ready_i_0_6[2] = ready_o_1_6[1];
    vc_i_0_6[0] = vc_i[0][6];
    data_i_0_6[0] = data_i[0][6];
    valid_i_0_6[0] = valid_i[0][6];
    ready_i_0_6[0] = ready_i[0][6];
end


/*Router 0,7*/    
cast_router #(
    .routing_table                  (routing_table_0_7)
)router_0_7(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_0_7),
    .data_i                         (data_i_0_7),
    .valid_i                        (valid_i_0_7),
    .ready_o                        (ready_o_0_7),
    .vc_o                           (vc_o_0_7),
    .data_o                         (data_o_0_7),
    .valid_o                        (valid_o_0_7),
    .ready_i                        (ready_i_0_7)
);


always_comb begin
    vc_i_0_7[3] = vc_o_0_6[4];
    data_i_0_7[3] = data_o_0_6[4];
    valid_i_0_7[3] = valid_o_0_6[4];
    ready_i_0_7[3] = ready_o_0_6[4];
    vc_i_0_7[2] = vc_o_1_7[1];
    data_i_0_7[2] = data_o_1_7[1];
    valid_i_0_7[2] = valid_o_1_7[1];
    ready_i_0_7[2] = ready_o_1_7[1];
    vc_i_0_7[0] = vc_i[0][7];
    data_i_0_7[0] = data_i[0][7];
    valid_i_0_7[0] = valid_i[0][7];
    ready_i_0_7[0] = ready_i[0][7];
end


/*Router 1,0*/    
cast_router #(
    .routing_table                  (routing_table_1_0)
)router_1_0(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_1_0),
    .data_i                         (data_i_1_0),
    .valid_i                        (valid_i_1_0),
    .ready_o                        (ready_o_1_0),
    .vc_o                           (vc_o_1_0),
    .data_o                         (data_o_1_0),
    .valid_o                        (valid_o_1_0),
    .ready_i                        (ready_i_1_0)
);


always_comb begin
    vc_i_1_0[4] = vc_o_1_1[3];
    data_i_1_0[4] = data_o_1_1[3];
    valid_i_1_0[4] = valid_o_1_1[3];
    ready_i_1_0[4] = ready_o_1_1[3];
    vc_i_1_0[1] = vc_o_0_0[2];
    data_i_1_0[1] = data_o_0_0[2];
    valid_i_1_0[1] = valid_o_0_0[2];
    ready_i_1_0[1] = ready_o_0_0[2];
    vc_i_1_0[2] = vc_o_2_0[1];
    data_i_1_0[2] = data_o_2_0[1];
    valid_i_1_0[2] = valid_o_2_0[1];
    ready_i_1_0[2] = ready_o_2_0[1];
    vc_i_1_0[0] = vc_i[1][0];
    data_i_1_0[0] = data_i[1][0];
    valid_i_1_0[0] = valid_i[1][0];
    ready_i_1_0[0] = ready_i[1][0];
end


/*Router 1,1*/    
cast_router #(
    .routing_table                  (routing_table_1_1)
)router_1_1(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_1_1),
    .data_i                         (data_i_1_1),
    .valid_i                        (valid_i_1_1),
    .ready_o                        (ready_o_1_1),
    .vc_o                           (vc_o_1_1),
    .data_o                         (data_o_1_1),
    .valid_o                        (valid_o_1_1),
    .ready_i                        (ready_i_1_1)
);


always_comb begin
    vc_i_1_1[3] = vc_o_1_0[4];
    data_i_1_1[3] = data_o_1_0[4];
    valid_i_1_1[3] = valid_o_1_0[4];
    ready_i_1_1[3] = ready_o_1_0[4];
    vc_i_1_1[4] = vc_o_1_2[3];
    data_i_1_1[4] = data_o_1_2[3];
    valid_i_1_1[4] = valid_o_1_2[3];
    ready_i_1_1[4] = ready_o_1_2[3];
    vc_i_1_1[1] = vc_o_0_1[2];
    data_i_1_1[1] = data_o_0_1[2];
    valid_i_1_1[1] = valid_o_0_1[2];
    ready_i_1_1[1] = ready_o_0_1[2];
    vc_i_1_1[2] = vc_o_2_1[1];
    data_i_1_1[2] = data_o_2_1[1];
    valid_i_1_1[2] = valid_o_2_1[1];
    ready_i_1_1[2] = ready_o_2_1[1];
    vc_i_1_1[0] = vc_i[1][1];
    data_i_1_1[0] = data_i[1][1];
    valid_i_1_1[0] = valid_i[1][1];
    ready_i_1_1[0] = ready_i[1][1];
end


/*Router 1,2*/    
cast_router #(
    .routing_table                  (routing_table_1_2)
)router_1_2(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_1_2),
    .data_i                         (data_i_1_2),
    .valid_i                        (valid_i_1_2),
    .ready_o                        (ready_o_1_2),
    .vc_o                           (vc_o_1_2),
    .data_o                         (data_o_1_2),
    .valid_o                        (valid_o_1_2),
    .ready_i                        (ready_i_1_2)
);


always_comb begin
    vc_i_1_2[3] = vc_o_1_1[4];
    data_i_1_2[3] = data_o_1_1[4];
    valid_i_1_2[3] = valid_o_1_1[4];
    ready_i_1_2[3] = ready_o_1_1[4];
    vc_i_1_2[4] = vc_o_1_3[3];
    data_i_1_2[4] = data_o_1_3[3];
    valid_i_1_2[4] = valid_o_1_3[3];
    ready_i_1_2[4] = ready_o_1_3[3];
    vc_i_1_2[1] = vc_o_0_2[2];
    data_i_1_2[1] = data_o_0_2[2];
    valid_i_1_2[1] = valid_o_0_2[2];
    ready_i_1_2[1] = ready_o_0_2[2];
    vc_i_1_2[2] = vc_o_2_2[1];
    data_i_1_2[2] = data_o_2_2[1];
    valid_i_1_2[2] = valid_o_2_2[1];
    ready_i_1_2[2] = ready_o_2_2[1];
    vc_i_1_2[0] = vc_i[1][2];
    data_i_1_2[0] = data_i[1][2];
    valid_i_1_2[0] = valid_i[1][2];
    ready_i_1_2[0] = ready_i[1][2];
end


/*Router 1,3*/    
cast_router #(
    .routing_table                  (routing_table_1_3)
)router_1_3(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_1_3),
    .data_i                         (data_i_1_3),
    .valid_i                        (valid_i_1_3),
    .ready_o                        (ready_o_1_3),
    .vc_o                           (vc_o_1_3),
    .data_o                         (data_o_1_3),
    .valid_o                        (valid_o_1_3),
    .ready_i                        (ready_i_1_3)
);


always_comb begin
    vc_i_1_3[3] = vc_o_1_2[4];
    data_i_1_3[3] = data_o_1_2[4];
    valid_i_1_3[3] = valid_o_1_2[4];
    ready_i_1_3[3] = ready_o_1_2[4];
    vc_i_1_3[4] = vc_o_1_4[3];
    data_i_1_3[4] = data_o_1_4[3];
    valid_i_1_3[4] = valid_o_1_4[3];
    ready_i_1_3[4] = ready_o_1_4[3];
    vc_i_1_3[1] = vc_o_0_3[2];
    data_i_1_3[1] = data_o_0_3[2];
    valid_i_1_3[1] = valid_o_0_3[2];
    ready_i_1_3[1] = ready_o_0_3[2];
    vc_i_1_3[2] = vc_o_2_3[1];
    data_i_1_3[2] = data_o_2_3[1];
    valid_i_1_3[2] = valid_o_2_3[1];
    ready_i_1_3[2] = ready_o_2_3[1];
    vc_i_1_3[0] = vc_i[1][3];
    data_i_1_3[0] = data_i[1][3];
    valid_i_1_3[0] = valid_i[1][3];
    ready_i_1_3[0] = ready_i[1][3];
end


/*Router 1,4*/    
cast_router #(
    .routing_table                  (routing_table_1_4)
)router_1_4(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_1_4),
    .data_i                         (data_i_1_4),
    .valid_i                        (valid_i_1_4),
    .ready_o                        (ready_o_1_4),
    .vc_o                           (vc_o_1_4),
    .data_o                         (data_o_1_4),
    .valid_o                        (valid_o_1_4),
    .ready_i                        (ready_i_1_4)
);


always_comb begin
    vc_i_1_4[3] = vc_o_1_3[4];
    data_i_1_4[3] = data_o_1_3[4];
    valid_i_1_4[3] = valid_o_1_3[4];
    ready_i_1_4[3] = ready_o_1_3[4];
    vc_i_1_4[4] = vc_o_1_5[3];
    data_i_1_4[4] = data_o_1_5[3];
    valid_i_1_4[4] = valid_o_1_5[3];
    ready_i_1_4[4] = ready_o_1_5[3];
    vc_i_1_4[1] = vc_o_0_4[2];
    data_i_1_4[1] = data_o_0_4[2];
    valid_i_1_4[1] = valid_o_0_4[2];
    ready_i_1_4[1] = ready_o_0_4[2];
    vc_i_1_4[2] = vc_o_2_4[1];
    data_i_1_4[2] = data_o_2_4[1];
    valid_i_1_4[2] = valid_o_2_4[1];
    ready_i_1_4[2] = ready_o_2_4[1];
    vc_i_1_4[0] = vc_i[1][4];
    data_i_1_4[0] = data_i[1][4];
    valid_i_1_4[0] = valid_i[1][4];
    ready_i_1_4[0] = ready_i[1][4];
end


/*Router 1,5*/    
cast_router #(
    .routing_table                  (routing_table_1_5)
)router_1_5(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_1_5),
    .data_i                         (data_i_1_5),
    .valid_i                        (valid_i_1_5),
    .ready_o                        (ready_o_1_5),
    .vc_o                           (vc_o_1_5),
    .data_o                         (data_o_1_5),
    .valid_o                        (valid_o_1_5),
    .ready_i                        (ready_i_1_5)
);


always_comb begin
    vc_i_1_5[3] = vc_o_1_4[4];
    data_i_1_5[3] = data_o_1_4[4];
    valid_i_1_5[3] = valid_o_1_4[4];
    ready_i_1_5[3] = ready_o_1_4[4];
    vc_i_1_5[4] = vc_o_1_6[3];
    data_i_1_5[4] = data_o_1_6[3];
    valid_i_1_5[4] = valid_o_1_6[3];
    ready_i_1_5[4] = ready_o_1_6[3];
    vc_i_1_5[1] = vc_o_0_5[2];
    data_i_1_5[1] = data_o_0_5[2];
    valid_i_1_5[1] = valid_o_0_5[2];
    ready_i_1_5[1] = ready_o_0_5[2];
    vc_i_1_5[2] = vc_o_2_5[1];
    data_i_1_5[2] = data_o_2_5[1];
    valid_i_1_5[2] = valid_o_2_5[1];
    ready_i_1_5[2] = ready_o_2_5[1];
    vc_i_1_5[0] = vc_i[1][5];
    data_i_1_5[0] = data_i[1][5];
    valid_i_1_5[0] = valid_i[1][5];
    ready_i_1_5[0] = ready_i[1][5];
end


/*Router 1,6*/    
cast_router #(
    .routing_table                  (routing_table_1_6)
)router_1_6(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_1_6),
    .data_i                         (data_i_1_6),
    .valid_i                        (valid_i_1_6),
    .ready_o                        (ready_o_1_6),
    .vc_o                           (vc_o_1_6),
    .data_o                         (data_o_1_6),
    .valid_o                        (valid_o_1_6),
    .ready_i                        (ready_i_1_6)
);


always_comb begin
    vc_i_1_6[3] = vc_o_1_5[4];
    data_i_1_6[3] = data_o_1_5[4];
    valid_i_1_6[3] = valid_o_1_5[4];
    ready_i_1_6[3] = ready_o_1_5[4];
    vc_i_1_6[4] = vc_o_1_7[3];
    data_i_1_6[4] = data_o_1_7[3];
    valid_i_1_6[4] = valid_o_1_7[3];
    ready_i_1_6[4] = ready_o_1_7[3];
    vc_i_1_6[1] = vc_o_0_6[2];
    data_i_1_6[1] = data_o_0_6[2];
    valid_i_1_6[1] = valid_o_0_6[2];
    ready_i_1_6[1] = ready_o_0_6[2];
    vc_i_1_6[2] = vc_o_2_6[1];
    data_i_1_6[2] = data_o_2_6[1];
    valid_i_1_6[2] = valid_o_2_6[1];
    ready_i_1_6[2] = ready_o_2_6[1];
    vc_i_1_6[0] = vc_i[1][6];
    data_i_1_6[0] = data_i[1][6];
    valid_i_1_6[0] = valid_i[1][6];
    ready_i_1_6[0] = ready_i[1][6];
end


/*Router 1,7*/    
cast_router #(
    .routing_table                  (routing_table_1_7)
)router_1_7(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_1_7),
    .data_i                         (data_i_1_7),
    .valid_i                        (valid_i_1_7),
    .ready_o                        (ready_o_1_7),
    .vc_o                           (vc_o_1_7),
    .data_o                         (data_o_1_7),
    .valid_o                        (valid_o_1_7),
    .ready_i                        (ready_i_1_7)
);


always_comb begin
    vc_i_1_7[3] = vc_o_1_6[4];
    data_i_1_7[3] = data_o_1_6[4];
    valid_i_1_7[3] = valid_o_1_6[4];
    ready_i_1_7[3] = ready_o_1_6[4];
    vc_i_1_7[1] = vc_o_0_7[2];
    data_i_1_7[1] = data_o_0_7[2];
    valid_i_1_7[1] = valid_o_0_7[2];
    ready_i_1_7[1] = ready_o_0_7[2];
    vc_i_1_7[2] = vc_o_2_7[1];
    data_i_1_7[2] = data_o_2_7[1];
    valid_i_1_7[2] = valid_o_2_7[1];
    ready_i_1_7[2] = ready_o_2_7[1];
    vc_i_1_7[0] = vc_i[1][7];
    data_i_1_7[0] = data_i[1][7];
    valid_i_1_7[0] = valid_i[1][7];
    ready_i_1_7[0] = ready_i[1][7];
end


/*Router 2,0*/    
cast_router #(
    .routing_table                  (routing_table_2_0)
)router_2_0(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_2_0),
    .data_i                         (data_i_2_0),
    .valid_i                        (valid_i_2_0),
    .ready_o                        (ready_o_2_0),
    .vc_o                           (vc_o_2_0),
    .data_o                         (data_o_2_0),
    .valid_o                        (valid_o_2_0),
    .ready_i                        (ready_i_2_0)
);


always_comb begin
    vc_i_2_0[4] = vc_o_2_1[3];
    data_i_2_0[4] = data_o_2_1[3];
    valid_i_2_0[4] = valid_o_2_1[3];
    ready_i_2_0[4] = ready_o_2_1[3];
    vc_i_2_0[1] = vc_o_1_0[2];
    data_i_2_0[1] = data_o_1_0[2];
    valid_i_2_0[1] = valid_o_1_0[2];
    ready_i_2_0[1] = ready_o_1_0[2];
    vc_i_2_0[2] = vc_o_3_0[1];
    data_i_2_0[2] = data_o_3_0[1];
    valid_i_2_0[2] = valid_o_3_0[1];
    ready_i_2_0[2] = ready_o_3_0[1];
    vc_i_2_0[0] = vc_i[2][0];
    data_i_2_0[0] = data_i[2][0];
    valid_i_2_0[0] = valid_i[2][0];
    ready_i_2_0[0] = ready_i[2][0];
end


/*Router 2,1*/    
cast_router #(
    .routing_table                  (routing_table_2_1)
)router_2_1(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_2_1),
    .data_i                         (data_i_2_1),
    .valid_i                        (valid_i_2_1),
    .ready_o                        (ready_o_2_1),
    .vc_o                           (vc_o_2_1),
    .data_o                         (data_o_2_1),
    .valid_o                        (valid_o_2_1),
    .ready_i                        (ready_i_2_1)
);


always_comb begin
    vc_i_2_1[3] = vc_o_2_0[4];
    data_i_2_1[3] = data_o_2_0[4];
    valid_i_2_1[3] = valid_o_2_0[4];
    ready_i_2_1[3] = ready_o_2_0[4];
    vc_i_2_1[4] = vc_o_2_2[3];
    data_i_2_1[4] = data_o_2_2[3];
    valid_i_2_1[4] = valid_o_2_2[3];
    ready_i_2_1[4] = ready_o_2_2[3];
    vc_i_2_1[1] = vc_o_1_1[2];
    data_i_2_1[1] = data_o_1_1[2];
    valid_i_2_1[1] = valid_o_1_1[2];
    ready_i_2_1[1] = ready_o_1_1[2];
    vc_i_2_1[2] = vc_o_3_1[1];
    data_i_2_1[2] = data_o_3_1[1];
    valid_i_2_1[2] = valid_o_3_1[1];
    ready_i_2_1[2] = ready_o_3_1[1];
    vc_i_2_1[0] = vc_i[2][1];
    data_i_2_1[0] = data_i[2][1];
    valid_i_2_1[0] = valid_i[2][1];
    ready_i_2_1[0] = ready_i[2][1];
end


/*Router 2,2*/    
cast_router #(
    .routing_table                  (routing_table_2_2)
)router_2_2(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_2_2),
    .data_i                         (data_i_2_2),
    .valid_i                        (valid_i_2_2),
    .ready_o                        (ready_o_2_2),
    .vc_o                           (vc_o_2_2),
    .data_o                         (data_o_2_2),
    .valid_o                        (valid_o_2_2),
    .ready_i                        (ready_i_2_2)
);


always_comb begin
    vc_i_2_2[3] = vc_o_2_1[4];
    data_i_2_2[3] = data_o_2_1[4];
    valid_i_2_2[3] = valid_o_2_1[4];
    ready_i_2_2[3] = ready_o_2_1[4];
    vc_i_2_2[4] = vc_o_2_3[3];
    data_i_2_2[4] = data_o_2_3[3];
    valid_i_2_2[4] = valid_o_2_3[3];
    ready_i_2_2[4] = ready_o_2_3[3];
    vc_i_2_2[1] = vc_o_1_2[2];
    data_i_2_2[1] = data_o_1_2[2];
    valid_i_2_2[1] = valid_o_1_2[2];
    ready_i_2_2[1] = ready_o_1_2[2];
    vc_i_2_2[2] = vc_o_3_2[1];
    data_i_2_2[2] = data_o_3_2[1];
    valid_i_2_2[2] = valid_o_3_2[1];
    ready_i_2_2[2] = ready_o_3_2[1];
    vc_i_2_2[0] = vc_i[2][2];
    data_i_2_2[0] = data_i[2][2];
    valid_i_2_2[0] = valid_i[2][2];
    ready_i_2_2[0] = ready_i[2][2];
end


/*Router 2,3*/    
cast_router #(
    .routing_table                  (routing_table_2_3)
)router_2_3(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_2_3),
    .data_i                         (data_i_2_3),
    .valid_i                        (valid_i_2_3),
    .ready_o                        (ready_o_2_3),
    .vc_o                           (vc_o_2_3),
    .data_o                         (data_o_2_3),
    .valid_o                        (valid_o_2_3),
    .ready_i                        (ready_i_2_3)
);


always_comb begin
    vc_i_2_3[3] = vc_o_2_2[4];
    data_i_2_3[3] = data_o_2_2[4];
    valid_i_2_3[3] = valid_o_2_2[4];
    ready_i_2_3[3] = ready_o_2_2[4];
    vc_i_2_3[4] = vc_o_2_4[3];
    data_i_2_3[4] = data_o_2_4[3];
    valid_i_2_3[4] = valid_o_2_4[3];
    ready_i_2_3[4] = ready_o_2_4[3];
    vc_i_2_3[1] = vc_o_1_3[2];
    data_i_2_3[1] = data_o_1_3[2];
    valid_i_2_3[1] = valid_o_1_3[2];
    ready_i_2_3[1] = ready_o_1_3[2];
    vc_i_2_3[2] = vc_o_3_3[1];
    data_i_2_3[2] = data_o_3_3[1];
    valid_i_2_3[2] = valid_o_3_3[1];
    ready_i_2_3[2] = ready_o_3_3[1];
    vc_i_2_3[0] = vc_i[2][3];
    data_i_2_3[0] = data_i[2][3];
    valid_i_2_3[0] = valid_i[2][3];
    ready_i_2_3[0] = ready_i[2][3];
end


/*Router 2,4*/    
cast_router #(
    .routing_table                  (routing_table_2_4)
)router_2_4(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_2_4),
    .data_i                         (data_i_2_4),
    .valid_i                        (valid_i_2_4),
    .ready_o                        (ready_o_2_4),
    .vc_o                           (vc_o_2_4),
    .data_o                         (data_o_2_4),
    .valid_o                        (valid_o_2_4),
    .ready_i                        (ready_i_2_4)
);


always_comb begin
    vc_i_2_4[3] = vc_o_2_3[4];
    data_i_2_4[3] = data_o_2_3[4];
    valid_i_2_4[3] = valid_o_2_3[4];
    ready_i_2_4[3] = ready_o_2_3[4];
    vc_i_2_4[4] = vc_o_2_5[3];
    data_i_2_4[4] = data_o_2_5[3];
    valid_i_2_4[4] = valid_o_2_5[3];
    ready_i_2_4[4] = ready_o_2_5[3];
    vc_i_2_4[1] = vc_o_1_4[2];
    data_i_2_4[1] = data_o_1_4[2];
    valid_i_2_4[1] = valid_o_1_4[2];
    ready_i_2_4[1] = ready_o_1_4[2];
    vc_i_2_4[2] = vc_o_3_4[1];
    data_i_2_4[2] = data_o_3_4[1];
    valid_i_2_4[2] = valid_o_3_4[1];
    ready_i_2_4[2] = ready_o_3_4[1];
    vc_i_2_4[0] = vc_i[2][4];
    data_i_2_4[0] = data_i[2][4];
    valid_i_2_4[0] = valid_i[2][4];
    ready_i_2_4[0] = ready_i[2][4];
end


/*Router 2,5*/    
cast_router #(
    .routing_table                  (routing_table_2_5)
)router_2_5(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_2_5),
    .data_i                         (data_i_2_5),
    .valid_i                        (valid_i_2_5),
    .ready_o                        (ready_o_2_5),
    .vc_o                           (vc_o_2_5),
    .data_o                         (data_o_2_5),
    .valid_o                        (valid_o_2_5),
    .ready_i                        (ready_i_2_5)
);


always_comb begin
    vc_i_2_5[3] = vc_o_2_4[4];
    data_i_2_5[3] = data_o_2_4[4];
    valid_i_2_5[3] = valid_o_2_4[4];
    ready_i_2_5[3] = ready_o_2_4[4];
    vc_i_2_5[4] = vc_o_2_6[3];
    data_i_2_5[4] = data_o_2_6[3];
    valid_i_2_5[4] = valid_o_2_6[3];
    ready_i_2_5[4] = ready_o_2_6[3];
    vc_i_2_5[1] = vc_o_1_5[2];
    data_i_2_5[1] = data_o_1_5[2];
    valid_i_2_5[1] = valid_o_1_5[2];
    ready_i_2_5[1] = ready_o_1_5[2];
    vc_i_2_5[2] = vc_o_3_5[1];
    data_i_2_5[2] = data_o_3_5[1];
    valid_i_2_5[2] = valid_o_3_5[1];
    ready_i_2_5[2] = ready_o_3_5[1];
    vc_i_2_5[0] = vc_i[2][5];
    data_i_2_5[0] = data_i[2][5];
    valid_i_2_5[0] = valid_i[2][5];
    ready_i_2_5[0] = ready_i[2][5];
end


/*Router 2,6*/    
cast_router #(
    .routing_table                  (routing_table_2_6)
)router_2_6(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_2_6),
    .data_i                         (data_i_2_6),
    .valid_i                        (valid_i_2_6),
    .ready_o                        (ready_o_2_6),
    .vc_o                           (vc_o_2_6),
    .data_o                         (data_o_2_6),
    .valid_o                        (valid_o_2_6),
    .ready_i                        (ready_i_2_6)
);


always_comb begin
    vc_i_2_6[3] = vc_o_2_5[4];
    data_i_2_6[3] = data_o_2_5[4];
    valid_i_2_6[3] = valid_o_2_5[4];
    ready_i_2_6[3] = ready_o_2_5[4];
    vc_i_2_6[4] = vc_o_2_7[3];
    data_i_2_6[4] = data_o_2_7[3];
    valid_i_2_6[4] = valid_o_2_7[3];
    ready_i_2_6[4] = ready_o_2_7[3];
    vc_i_2_6[1] = vc_o_1_6[2];
    data_i_2_6[1] = data_o_1_6[2];
    valid_i_2_6[1] = valid_o_1_6[2];
    ready_i_2_6[1] = ready_o_1_6[2];
    vc_i_2_6[2] = vc_o_3_6[1];
    data_i_2_6[2] = data_o_3_6[1];
    valid_i_2_6[2] = valid_o_3_6[1];
    ready_i_2_6[2] = ready_o_3_6[1];
    vc_i_2_6[0] = vc_i[2][6];
    data_i_2_6[0] = data_i[2][6];
    valid_i_2_6[0] = valid_i[2][6];
    ready_i_2_6[0] = ready_i[2][6];
end


/*Router 2,7*/    
cast_router #(
    .routing_table                  (routing_table_2_7)
)router_2_7(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_2_7),
    .data_i                         (data_i_2_7),
    .valid_i                        (valid_i_2_7),
    .ready_o                        (ready_o_2_7),
    .vc_o                           (vc_o_2_7),
    .data_o                         (data_o_2_7),
    .valid_o                        (valid_o_2_7),
    .ready_i                        (ready_i_2_7)
);


always_comb begin
    vc_i_2_7[3] = vc_o_2_6[4];
    data_i_2_7[3] = data_o_2_6[4];
    valid_i_2_7[3] = valid_o_2_6[4];
    ready_i_2_7[3] = ready_o_2_6[4];
    vc_i_2_7[1] = vc_o_1_7[2];
    data_i_2_7[1] = data_o_1_7[2];
    valid_i_2_7[1] = valid_o_1_7[2];
    ready_i_2_7[1] = ready_o_1_7[2];
    vc_i_2_7[2] = vc_o_3_7[1];
    data_i_2_7[2] = data_o_3_7[1];
    valid_i_2_7[2] = valid_o_3_7[1];
    ready_i_2_7[2] = ready_o_3_7[1];
    vc_i_2_7[0] = vc_i[2][7];
    data_i_2_7[0] = data_i[2][7];
    valid_i_2_7[0] = valid_i[2][7];
    ready_i_2_7[0] = ready_i[2][7];
end


/*Router 3,0*/    
cast_router #(
    .routing_table                  (routing_table_3_0)
)router_3_0(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_3_0),
    .data_i                         (data_i_3_0),
    .valid_i                        (valid_i_3_0),
    .ready_o                        (ready_o_3_0),
    .vc_o                           (vc_o_3_0),
    .data_o                         (data_o_3_0),
    .valid_o                        (valid_o_3_0),
    .ready_i                        (ready_i_3_0)
);


always_comb begin
    vc_i_3_0[4] = vc_o_3_1[3];
    data_i_3_0[4] = data_o_3_1[3];
    valid_i_3_0[4] = valid_o_3_1[3];
    ready_i_3_0[4] = ready_o_3_1[3];
    vc_i_3_0[1] = vc_o_2_0[2];
    data_i_3_0[1] = data_o_2_0[2];
    valid_i_3_0[1] = valid_o_2_0[2];
    ready_i_3_0[1] = ready_o_2_0[2];
    vc_i_3_0[2] = vc_o_4_0[1];
    data_i_3_0[2] = data_o_4_0[1];
    valid_i_3_0[2] = valid_o_4_0[1];
    ready_i_3_0[2] = ready_o_4_0[1];
    vc_i_3_0[0] = vc_i[3][0];
    data_i_3_0[0] = data_i[3][0];
    valid_i_3_0[0] = valid_i[3][0];
    ready_i_3_0[0] = ready_i[3][0];
end


/*Router 3,1*/    
cast_router #(
    .routing_table                  (routing_table_3_1)
)router_3_1(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_3_1),
    .data_i                         (data_i_3_1),
    .valid_i                        (valid_i_3_1),
    .ready_o                        (ready_o_3_1),
    .vc_o                           (vc_o_3_1),
    .data_o                         (data_o_3_1),
    .valid_o                        (valid_o_3_1),
    .ready_i                        (ready_i_3_1)
);


always_comb begin
    vc_i_3_1[3] = vc_o_3_0[4];
    data_i_3_1[3] = data_o_3_0[4];
    valid_i_3_1[3] = valid_o_3_0[4];
    ready_i_3_1[3] = ready_o_3_0[4];
    vc_i_3_1[4] = vc_o_3_2[3];
    data_i_3_1[4] = data_o_3_2[3];
    valid_i_3_1[4] = valid_o_3_2[3];
    ready_i_3_1[4] = ready_o_3_2[3];
    vc_i_3_1[1] = vc_o_2_1[2];
    data_i_3_1[1] = data_o_2_1[2];
    valid_i_3_1[1] = valid_o_2_1[2];
    ready_i_3_1[1] = ready_o_2_1[2];
    vc_i_3_1[2] = vc_o_4_1[1];
    data_i_3_1[2] = data_o_4_1[1];
    valid_i_3_1[2] = valid_o_4_1[1];
    ready_i_3_1[2] = ready_o_4_1[1];
    vc_i_3_1[0] = vc_i[3][1];
    data_i_3_1[0] = data_i[3][1];
    valid_i_3_1[0] = valid_i[3][1];
    ready_i_3_1[0] = ready_i[3][1];
end


/*Router 3,2*/    
cast_router #(
    .routing_table                  (routing_table_3_2)
)router_3_2(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_3_2),
    .data_i                         (data_i_3_2),
    .valid_i                        (valid_i_3_2),
    .ready_o                        (ready_o_3_2),
    .vc_o                           (vc_o_3_2),
    .data_o                         (data_o_3_2),
    .valid_o                        (valid_o_3_2),
    .ready_i                        (ready_i_3_2)
);


always_comb begin
    vc_i_3_2[3] = vc_o_3_1[4];
    data_i_3_2[3] = data_o_3_1[4];
    valid_i_3_2[3] = valid_o_3_1[4];
    ready_i_3_2[3] = ready_o_3_1[4];
    vc_i_3_2[4] = vc_o_3_3[3];
    data_i_3_2[4] = data_o_3_3[3];
    valid_i_3_2[4] = valid_o_3_3[3];
    ready_i_3_2[4] = ready_o_3_3[3];
    vc_i_3_2[1] = vc_o_2_2[2];
    data_i_3_2[1] = data_o_2_2[2];
    valid_i_3_2[1] = valid_o_2_2[2];
    ready_i_3_2[1] = ready_o_2_2[2];
    vc_i_3_2[2] = vc_o_4_2[1];
    data_i_3_2[2] = data_o_4_2[1];
    valid_i_3_2[2] = valid_o_4_2[1];
    ready_i_3_2[2] = ready_o_4_2[1];
    vc_i_3_2[0] = vc_i[3][2];
    data_i_3_2[0] = data_i[3][2];
    valid_i_3_2[0] = valid_i[3][2];
    ready_i_3_2[0] = ready_i[3][2];
end


/*Router 3,3*/    
cast_router #(
    .routing_table                  (routing_table_3_3)
)router_3_3(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_3_3),
    .data_i                         (data_i_3_3),
    .valid_i                        (valid_i_3_3),
    .ready_o                        (ready_o_3_3),
    .vc_o                           (vc_o_3_3),
    .data_o                         (data_o_3_3),
    .valid_o                        (valid_o_3_3),
    .ready_i                        (ready_i_3_3)
);


always_comb begin
    vc_i_3_3[3] = vc_o_3_2[4];
    data_i_3_3[3] = data_o_3_2[4];
    valid_i_3_3[3] = valid_o_3_2[4];
    ready_i_3_3[3] = ready_o_3_2[4];
    vc_i_3_3[4] = vc_o_3_4[3];
    data_i_3_3[4] = data_o_3_4[3];
    valid_i_3_3[4] = valid_o_3_4[3];
    ready_i_3_3[4] = ready_o_3_4[3];
    vc_i_3_3[1] = vc_o_2_3[2];
    data_i_3_3[1] = data_o_2_3[2];
    valid_i_3_3[1] = valid_o_2_3[2];
    ready_i_3_3[1] = ready_o_2_3[2];
    vc_i_3_3[2] = vc_o_4_3[1];
    data_i_3_3[2] = data_o_4_3[1];
    valid_i_3_3[2] = valid_o_4_3[1];
    ready_i_3_3[2] = ready_o_4_3[1];
    vc_i_3_3[0] = vc_i[3][3];
    data_i_3_3[0] = data_i[3][3];
    valid_i_3_3[0] = valid_i[3][3];
    ready_i_3_3[0] = ready_i[3][3];
end


/*Router 3,4*/    
cast_router #(
    .routing_table                  (routing_table_3_4)
)router_3_4(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_3_4),
    .data_i                         (data_i_3_4),
    .valid_i                        (valid_i_3_4),
    .ready_o                        (ready_o_3_4),
    .vc_o                           (vc_o_3_4),
    .data_o                         (data_o_3_4),
    .valid_o                        (valid_o_3_4),
    .ready_i                        (ready_i_3_4)
);


always_comb begin
    vc_i_3_4[3] = vc_o_3_3[4];
    data_i_3_4[3] = data_o_3_3[4];
    valid_i_3_4[3] = valid_o_3_3[4];
    ready_i_3_4[3] = ready_o_3_3[4];
    vc_i_3_4[4] = vc_o_3_5[3];
    data_i_3_4[4] = data_o_3_5[3];
    valid_i_3_4[4] = valid_o_3_5[3];
    ready_i_3_4[4] = ready_o_3_5[3];
    vc_i_3_4[1] = vc_o_2_4[2];
    data_i_3_4[1] = data_o_2_4[2];
    valid_i_3_4[1] = valid_o_2_4[2];
    ready_i_3_4[1] = ready_o_2_4[2];
    vc_i_3_4[2] = vc_o_4_4[1];
    data_i_3_4[2] = data_o_4_4[1];
    valid_i_3_4[2] = valid_o_4_4[1];
    ready_i_3_4[2] = ready_o_4_4[1];
    vc_i_3_4[0] = vc_i[3][4];
    data_i_3_4[0] = data_i[3][4];
    valid_i_3_4[0] = valid_i[3][4];
    ready_i_3_4[0] = ready_i[3][4];
end


/*Router 3,5*/    
cast_router #(
    .routing_table                  (routing_table_3_5)
)router_3_5(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_3_5),
    .data_i                         (data_i_3_5),
    .valid_i                        (valid_i_3_5),
    .ready_o                        (ready_o_3_5),
    .vc_o                           (vc_o_3_5),
    .data_o                         (data_o_3_5),
    .valid_o                        (valid_o_3_5),
    .ready_i                        (ready_i_3_5)
);


always_comb begin
    vc_i_3_5[3] = vc_o_3_4[4];
    data_i_3_5[3] = data_o_3_4[4];
    valid_i_3_5[3] = valid_o_3_4[4];
    ready_i_3_5[3] = ready_o_3_4[4];
    vc_i_3_5[4] = vc_o_3_6[3];
    data_i_3_5[4] = data_o_3_6[3];
    valid_i_3_5[4] = valid_o_3_6[3];
    ready_i_3_5[4] = ready_o_3_6[3];
    vc_i_3_5[1] = vc_o_2_5[2];
    data_i_3_5[1] = data_o_2_5[2];
    valid_i_3_5[1] = valid_o_2_5[2];
    ready_i_3_5[1] = ready_o_2_5[2];
    vc_i_3_5[2] = vc_o_4_5[1];
    data_i_3_5[2] = data_o_4_5[1];
    valid_i_3_5[2] = valid_o_4_5[1];
    ready_i_3_5[2] = ready_o_4_5[1];
    vc_i_3_5[0] = vc_i[3][5];
    data_i_3_5[0] = data_i[3][5];
    valid_i_3_5[0] = valid_i[3][5];
    ready_i_3_5[0] = ready_i[3][5];
end


/*Router 3,6*/    
cast_router #(
    .routing_table                  (routing_table_3_6)
)router_3_6(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_3_6),
    .data_i                         (data_i_3_6),
    .valid_i                        (valid_i_3_6),
    .ready_o                        (ready_o_3_6),
    .vc_o                           (vc_o_3_6),
    .data_o                         (data_o_3_6),
    .valid_o                        (valid_o_3_6),
    .ready_i                        (ready_i_3_6)
);


always_comb begin
    vc_i_3_6[3] = vc_o_3_5[4];
    data_i_3_6[3] = data_o_3_5[4];
    valid_i_3_6[3] = valid_o_3_5[4];
    ready_i_3_6[3] = ready_o_3_5[4];
    vc_i_3_6[4] = vc_o_3_7[3];
    data_i_3_6[4] = data_o_3_7[3];
    valid_i_3_6[4] = valid_o_3_7[3];
    ready_i_3_6[4] = ready_o_3_7[3];
    vc_i_3_6[1] = vc_o_2_6[2];
    data_i_3_6[1] = data_o_2_6[2];
    valid_i_3_6[1] = valid_o_2_6[2];
    ready_i_3_6[1] = ready_o_2_6[2];
    vc_i_3_6[2] = vc_o_4_6[1];
    data_i_3_6[2] = data_o_4_6[1];
    valid_i_3_6[2] = valid_o_4_6[1];
    ready_i_3_6[2] = ready_o_4_6[1];
    vc_i_3_6[0] = vc_i[3][6];
    data_i_3_6[0] = data_i[3][6];
    valid_i_3_6[0] = valid_i[3][6];
    ready_i_3_6[0] = ready_i[3][6];
end


/*Router 3,7*/    
cast_router #(
    .routing_table                  (routing_table_3_7)
)router_3_7(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_3_7),
    .data_i                         (data_i_3_7),
    .valid_i                        (valid_i_3_7),
    .ready_o                        (ready_o_3_7),
    .vc_o                           (vc_o_3_7),
    .data_o                         (data_o_3_7),
    .valid_o                        (valid_o_3_7),
    .ready_i                        (ready_i_3_7)
);


always_comb begin
    vc_i_3_7[3] = vc_o_3_6[4];
    data_i_3_7[3] = data_o_3_6[4];
    valid_i_3_7[3] = valid_o_3_6[4];
    ready_i_3_7[3] = ready_o_3_6[4];
    vc_i_3_7[1] = vc_o_2_7[2];
    data_i_3_7[1] = data_o_2_7[2];
    valid_i_3_7[1] = valid_o_2_7[2];
    ready_i_3_7[1] = ready_o_2_7[2];
    vc_i_3_7[2] = vc_o_4_7[1];
    data_i_3_7[2] = data_o_4_7[1];
    valid_i_3_7[2] = valid_o_4_7[1];
    ready_i_3_7[2] = ready_o_4_7[1];
    vc_i_3_7[0] = vc_i[3][7];
    data_i_3_7[0] = data_i[3][7];
    valid_i_3_7[0] = valid_i[3][7];
    ready_i_3_7[0] = ready_i[3][7];
end


/*Router 4,0*/    
cast_router #(
    .routing_table                  (routing_table_4_0)
)router_4_0(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_4_0),
    .data_i                         (data_i_4_0),
    .valid_i                        (valid_i_4_0),
    .ready_o                        (ready_o_4_0),
    .vc_o                           (vc_o_4_0),
    .data_o                         (data_o_4_0),
    .valid_o                        (valid_o_4_0),
    .ready_i                        (ready_i_4_0)
);


always_comb begin
    vc_i_4_0[4] = vc_o_4_1[3];
    data_i_4_0[4] = data_o_4_1[3];
    valid_i_4_0[4] = valid_o_4_1[3];
    ready_i_4_0[4] = ready_o_4_1[3];
    vc_i_4_0[1] = vc_o_3_0[2];
    data_i_4_0[1] = data_o_3_0[2];
    valid_i_4_0[1] = valid_o_3_0[2];
    ready_i_4_0[1] = ready_o_3_0[2];
    vc_i_4_0[2] = vc_o_5_0[1];
    data_i_4_0[2] = data_o_5_0[1];
    valid_i_4_0[2] = valid_o_5_0[1];
    ready_i_4_0[2] = ready_o_5_0[1];
    vc_i_4_0[0] = vc_i[4][0];
    data_i_4_0[0] = data_i[4][0];
    valid_i_4_0[0] = valid_i[4][0];
    ready_i_4_0[0] = ready_i[4][0];
end


/*Router 4,1*/    
cast_router #(
    .routing_table                  (routing_table_4_1)
)router_4_1(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_4_1),
    .data_i                         (data_i_4_1),
    .valid_i                        (valid_i_4_1),
    .ready_o                        (ready_o_4_1),
    .vc_o                           (vc_o_4_1),
    .data_o                         (data_o_4_1),
    .valid_o                        (valid_o_4_1),
    .ready_i                        (ready_i_4_1)
);


always_comb begin
    vc_i_4_1[3] = vc_o_4_0[4];
    data_i_4_1[3] = data_o_4_0[4];
    valid_i_4_1[3] = valid_o_4_0[4];
    ready_i_4_1[3] = ready_o_4_0[4];
    vc_i_4_1[4] = vc_o_4_2[3];
    data_i_4_1[4] = data_o_4_2[3];
    valid_i_4_1[4] = valid_o_4_2[3];
    ready_i_4_1[4] = ready_o_4_2[3];
    vc_i_4_1[1] = vc_o_3_1[2];
    data_i_4_1[1] = data_o_3_1[2];
    valid_i_4_1[1] = valid_o_3_1[2];
    ready_i_4_1[1] = ready_o_3_1[2];
    vc_i_4_1[2] = vc_o_5_1[1];
    data_i_4_1[2] = data_o_5_1[1];
    valid_i_4_1[2] = valid_o_5_1[1];
    ready_i_4_1[2] = ready_o_5_1[1];
    vc_i_4_1[0] = vc_i[4][1];
    data_i_4_1[0] = data_i[4][1];
    valid_i_4_1[0] = valid_i[4][1];
    ready_i_4_1[0] = ready_i[4][1];
end


/*Router 4,2*/    
cast_router #(
    .routing_table                  (routing_table_4_2)
)router_4_2(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_4_2),
    .data_i                         (data_i_4_2),
    .valid_i                        (valid_i_4_2),
    .ready_o                        (ready_o_4_2),
    .vc_o                           (vc_o_4_2),
    .data_o                         (data_o_4_2),
    .valid_o                        (valid_o_4_2),
    .ready_i                        (ready_i_4_2)
);


always_comb begin
    vc_i_4_2[3] = vc_o_4_1[4];
    data_i_4_2[3] = data_o_4_1[4];
    valid_i_4_2[3] = valid_o_4_1[4];
    ready_i_4_2[3] = ready_o_4_1[4];
    vc_i_4_2[4] = vc_o_4_3[3];
    data_i_4_2[4] = data_o_4_3[3];
    valid_i_4_2[4] = valid_o_4_3[3];
    ready_i_4_2[4] = ready_o_4_3[3];
    vc_i_4_2[1] = vc_o_3_2[2];
    data_i_4_2[1] = data_o_3_2[2];
    valid_i_4_2[1] = valid_o_3_2[2];
    ready_i_4_2[1] = ready_o_3_2[2];
    vc_i_4_2[2] = vc_o_5_2[1];
    data_i_4_2[2] = data_o_5_2[1];
    valid_i_4_2[2] = valid_o_5_2[1];
    ready_i_4_2[2] = ready_o_5_2[1];
    vc_i_4_2[0] = vc_i[4][2];
    data_i_4_2[0] = data_i[4][2];
    valid_i_4_2[0] = valid_i[4][2];
    ready_i_4_2[0] = ready_i[4][2];
end


/*Router 4,3*/    
cast_router #(
    .routing_table                  (routing_table_4_3)
)router_4_3(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_4_3),
    .data_i                         (data_i_4_3),
    .valid_i                        (valid_i_4_3),
    .ready_o                        (ready_o_4_3),
    .vc_o                           (vc_o_4_3),
    .data_o                         (data_o_4_3),
    .valid_o                        (valid_o_4_3),
    .ready_i                        (ready_i_4_3)
);


always_comb begin
    vc_i_4_3[3] = vc_o_4_2[4];
    data_i_4_3[3] = data_o_4_2[4];
    valid_i_4_3[3] = valid_o_4_2[4];
    ready_i_4_3[3] = ready_o_4_2[4];
    vc_i_4_3[4] = vc_o_4_4[3];
    data_i_4_3[4] = data_o_4_4[3];
    valid_i_4_3[4] = valid_o_4_4[3];
    ready_i_4_3[4] = ready_o_4_4[3];
    vc_i_4_3[1] = vc_o_3_3[2];
    data_i_4_3[1] = data_o_3_3[2];
    valid_i_4_3[1] = valid_o_3_3[2];
    ready_i_4_3[1] = ready_o_3_3[2];
    vc_i_4_3[2] = vc_o_5_3[1];
    data_i_4_3[2] = data_o_5_3[1];
    valid_i_4_3[2] = valid_o_5_3[1];
    ready_i_4_3[2] = ready_o_5_3[1];
    vc_i_4_3[0] = vc_i[4][3];
    data_i_4_3[0] = data_i[4][3];
    valid_i_4_3[0] = valid_i[4][3];
    ready_i_4_3[0] = ready_i[4][3];
end


/*Router 4,4*/    
cast_router #(
    .routing_table                  (routing_table_4_4)
)router_4_4(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_4_4),
    .data_i                         (data_i_4_4),
    .valid_i                        (valid_i_4_4),
    .ready_o                        (ready_o_4_4),
    .vc_o                           (vc_o_4_4),
    .data_o                         (data_o_4_4),
    .valid_o                        (valid_o_4_4),
    .ready_i                        (ready_i_4_4)
);


always_comb begin
    vc_i_4_4[3] = vc_o_4_3[4];
    data_i_4_4[3] = data_o_4_3[4];
    valid_i_4_4[3] = valid_o_4_3[4];
    ready_i_4_4[3] = ready_o_4_3[4];
    vc_i_4_4[4] = vc_o_4_5[3];
    data_i_4_4[4] = data_o_4_5[3];
    valid_i_4_4[4] = valid_o_4_5[3];
    ready_i_4_4[4] = ready_o_4_5[3];
    vc_i_4_4[1] = vc_o_3_4[2];
    data_i_4_4[1] = data_o_3_4[2];
    valid_i_4_4[1] = valid_o_3_4[2];
    ready_i_4_4[1] = ready_o_3_4[2];
    vc_i_4_4[2] = vc_o_5_4[1];
    data_i_4_4[2] = data_o_5_4[1];
    valid_i_4_4[2] = valid_o_5_4[1];
    ready_i_4_4[2] = ready_o_5_4[1];
    vc_i_4_4[0] = vc_i[4][4];
    data_i_4_4[0] = data_i[4][4];
    valid_i_4_4[0] = valid_i[4][4];
    ready_i_4_4[0] = ready_i[4][4];
end


/*Router 4,5*/    
cast_router #(
    .routing_table                  (routing_table_4_5)
)router_4_5(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_4_5),
    .data_i                         (data_i_4_5),
    .valid_i                        (valid_i_4_5),
    .ready_o                        (ready_o_4_5),
    .vc_o                           (vc_o_4_5),
    .data_o                         (data_o_4_5),
    .valid_o                        (valid_o_4_5),
    .ready_i                        (ready_i_4_5)
);


always_comb begin
    vc_i_4_5[3] = vc_o_4_4[4];
    data_i_4_5[3] = data_o_4_4[4];
    valid_i_4_5[3] = valid_o_4_4[4];
    ready_i_4_5[3] = ready_o_4_4[4];
    vc_i_4_5[4] = vc_o_4_6[3];
    data_i_4_5[4] = data_o_4_6[3];
    valid_i_4_5[4] = valid_o_4_6[3];
    ready_i_4_5[4] = ready_o_4_6[3];
    vc_i_4_5[1] = vc_o_3_5[2];
    data_i_4_5[1] = data_o_3_5[2];
    valid_i_4_5[1] = valid_o_3_5[2];
    ready_i_4_5[1] = ready_o_3_5[2];
    vc_i_4_5[2] = vc_o_5_5[1];
    data_i_4_5[2] = data_o_5_5[1];
    valid_i_4_5[2] = valid_o_5_5[1];
    ready_i_4_5[2] = ready_o_5_5[1];
    vc_i_4_5[0] = vc_i[4][5];
    data_i_4_5[0] = data_i[4][5];
    valid_i_4_5[0] = valid_i[4][5];
    ready_i_4_5[0] = ready_i[4][5];
end


/*Router 4,6*/    
cast_router #(
    .routing_table                  (routing_table_4_6)
)router_4_6(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_4_6),
    .data_i                         (data_i_4_6),
    .valid_i                        (valid_i_4_6),
    .ready_o                        (ready_o_4_6),
    .vc_o                           (vc_o_4_6),
    .data_o                         (data_o_4_6),
    .valid_o                        (valid_o_4_6),
    .ready_i                        (ready_i_4_6)
);


always_comb begin
    vc_i_4_6[3] = vc_o_4_5[4];
    data_i_4_6[3] = data_o_4_5[4];
    valid_i_4_6[3] = valid_o_4_5[4];
    ready_i_4_6[3] = ready_o_4_5[4];
    vc_i_4_6[4] = vc_o_4_7[3];
    data_i_4_6[4] = data_o_4_7[3];
    valid_i_4_6[4] = valid_o_4_7[3];
    ready_i_4_6[4] = ready_o_4_7[3];
    vc_i_4_6[1] = vc_o_3_6[2];
    data_i_4_6[1] = data_o_3_6[2];
    valid_i_4_6[1] = valid_o_3_6[2];
    ready_i_4_6[1] = ready_o_3_6[2];
    vc_i_4_6[2] = vc_o_5_6[1];
    data_i_4_6[2] = data_o_5_6[1];
    valid_i_4_6[2] = valid_o_5_6[1];
    ready_i_4_6[2] = ready_o_5_6[1];
    vc_i_4_6[0] = vc_i[4][6];
    data_i_4_6[0] = data_i[4][6];
    valid_i_4_6[0] = valid_i[4][6];
    ready_i_4_6[0] = ready_i[4][6];
end


/*Router 4,7*/    
cast_router #(
    .routing_table                  (routing_table_4_7)
)router_4_7(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_4_7),
    .data_i                         (data_i_4_7),
    .valid_i                        (valid_i_4_7),
    .ready_o                        (ready_o_4_7),
    .vc_o                           (vc_o_4_7),
    .data_o                         (data_o_4_7),
    .valid_o                        (valid_o_4_7),
    .ready_i                        (ready_i_4_7)
);


always_comb begin
    vc_i_4_7[3] = vc_o_4_6[4];
    data_i_4_7[3] = data_o_4_6[4];
    valid_i_4_7[3] = valid_o_4_6[4];
    ready_i_4_7[3] = ready_o_4_6[4];
    vc_i_4_7[1] = vc_o_3_7[2];
    data_i_4_7[1] = data_o_3_7[2];
    valid_i_4_7[1] = valid_o_3_7[2];
    ready_i_4_7[1] = ready_o_3_7[2];
    vc_i_4_7[2] = vc_o_5_7[1];
    data_i_4_7[2] = data_o_5_7[1];
    valid_i_4_7[2] = valid_o_5_7[1];
    ready_i_4_7[2] = ready_o_5_7[1];
    vc_i_4_7[0] = vc_i[4][7];
    data_i_4_7[0] = data_i[4][7];
    valid_i_4_7[0] = valid_i[4][7];
    ready_i_4_7[0] = ready_i[4][7];
end


/*Router 5,0*/    
cast_router #(
    .routing_table                  (routing_table_5_0)
)router_5_0(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_5_0),
    .data_i                         (data_i_5_0),
    .valid_i                        (valid_i_5_0),
    .ready_o                        (ready_o_5_0),
    .vc_o                           (vc_o_5_0),
    .data_o                         (data_o_5_0),
    .valid_o                        (valid_o_5_0),
    .ready_i                        (ready_i_5_0)
);


always_comb begin
    vc_i_5_0[4] = vc_o_5_1[3];
    data_i_5_0[4] = data_o_5_1[3];
    valid_i_5_0[4] = valid_o_5_1[3];
    ready_i_5_0[4] = ready_o_5_1[3];
    vc_i_5_0[1] = vc_o_4_0[2];
    data_i_5_0[1] = data_o_4_0[2];
    valid_i_5_0[1] = valid_o_4_0[2];
    ready_i_5_0[1] = ready_o_4_0[2];
    vc_i_5_0[0] = vc_i[5][0];
    data_i_5_0[0] = data_i[5][0];
    valid_i_5_0[0] = valid_i[5][0];
    ready_i_5_0[0] = ready_i[5][0];
end


/*Router 5,1*/    
cast_router #(
    .routing_table                  (routing_table_5_1)
)router_5_1(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_5_1),
    .data_i                         (data_i_5_1),
    .valid_i                        (valid_i_5_1),
    .ready_o                        (ready_o_5_1),
    .vc_o                           (vc_o_5_1),
    .data_o                         (data_o_5_1),
    .valid_o                        (valid_o_5_1),
    .ready_i                        (ready_i_5_1)
);


always_comb begin
    vc_i_5_1[3] = vc_o_5_0[4];
    data_i_5_1[3] = data_o_5_0[4];
    valid_i_5_1[3] = valid_o_5_0[4];
    ready_i_5_1[3] = ready_o_5_0[4];
    vc_i_5_1[4] = vc_o_5_2[3];
    data_i_5_1[4] = data_o_5_2[3];
    valid_i_5_1[4] = valid_o_5_2[3];
    ready_i_5_1[4] = ready_o_5_2[3];
    vc_i_5_1[1] = vc_o_4_1[2];
    data_i_5_1[1] = data_o_4_1[2];
    valid_i_5_1[1] = valid_o_4_1[2];
    ready_i_5_1[1] = ready_o_4_1[2];
    vc_i_5_1[0] = vc_i[5][1];
    data_i_5_1[0] = data_i[5][1];
    valid_i_5_1[0] = valid_i[5][1];
    ready_i_5_1[0] = ready_i[5][1];
end


/*Router 5,2*/    
cast_router #(
    .routing_table                  (routing_table_5_2)
)router_5_2(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_5_2),
    .data_i                         (data_i_5_2),
    .valid_i                        (valid_i_5_2),
    .ready_o                        (ready_o_5_2),
    .vc_o                           (vc_o_5_2),
    .data_o                         (data_o_5_2),
    .valid_o                        (valid_o_5_2),
    .ready_i                        (ready_i_5_2)
);


always_comb begin
    vc_i_5_2[3] = vc_o_5_1[4];
    data_i_5_2[3] = data_o_5_1[4];
    valid_i_5_2[3] = valid_o_5_1[4];
    ready_i_5_2[3] = ready_o_5_1[4];
    vc_i_5_2[4] = vc_o_5_3[3];
    data_i_5_2[4] = data_o_5_3[3];
    valid_i_5_2[4] = valid_o_5_3[3];
    ready_i_5_2[4] = ready_o_5_3[3];
    vc_i_5_2[1] = vc_o_4_2[2];
    data_i_5_2[1] = data_o_4_2[2];
    valid_i_5_2[1] = valid_o_4_2[2];
    ready_i_5_2[1] = ready_o_4_2[2];
    vc_i_5_2[0] = vc_i[5][2];
    data_i_5_2[0] = data_i[5][2];
    valid_i_5_2[0] = valid_i[5][2];
    ready_i_5_2[0] = ready_i[5][2];
end


/*Router 5,3*/    
cast_router #(
    .routing_table                  (routing_table_5_3)
)router_5_3(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_5_3),
    .data_i                         (data_i_5_3),
    .valid_i                        (valid_i_5_3),
    .ready_o                        (ready_o_5_3),
    .vc_o                           (vc_o_5_3),
    .data_o                         (data_o_5_3),
    .valid_o                        (valid_o_5_3),
    .ready_i                        (ready_i_5_3)
);


always_comb begin
    vc_i_5_3[3] = vc_o_5_2[4];
    data_i_5_3[3] = data_o_5_2[4];
    valid_i_5_3[3] = valid_o_5_2[4];
    ready_i_5_3[3] = ready_o_5_2[4];
    vc_i_5_3[4] = vc_o_5_4[3];
    data_i_5_3[4] = data_o_5_4[3];
    valid_i_5_3[4] = valid_o_5_4[3];
    ready_i_5_3[4] = ready_o_5_4[3];
    vc_i_5_3[1] = vc_o_4_3[2];
    data_i_5_3[1] = data_o_4_3[2];
    valid_i_5_3[1] = valid_o_4_3[2];
    ready_i_5_3[1] = ready_o_4_3[2];
    vc_i_5_3[0] = vc_i[5][3];
    data_i_5_3[0] = data_i[5][3];
    valid_i_5_3[0] = valid_i[5][3];
    ready_i_5_3[0] = ready_i[5][3];
end


/*Router 5,4*/    
cast_router #(
    .routing_table                  (routing_table_5_4)
)router_5_4(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_5_4),
    .data_i                         (data_i_5_4),
    .valid_i                        (valid_i_5_4),
    .ready_o                        (ready_o_5_4),
    .vc_o                           (vc_o_5_4),
    .data_o                         (data_o_5_4),
    .valid_o                        (valid_o_5_4),
    .ready_i                        (ready_i_5_4)
);


always_comb begin
    vc_i_5_4[3] = vc_o_5_3[4];
    data_i_5_4[3] = data_o_5_3[4];
    valid_i_5_4[3] = valid_o_5_3[4];
    ready_i_5_4[3] = ready_o_5_3[4];
    vc_i_5_4[4] = vc_o_5_5[3];
    data_i_5_4[4] = data_o_5_5[3];
    valid_i_5_4[4] = valid_o_5_5[3];
    ready_i_5_4[4] = ready_o_5_5[3];
    vc_i_5_4[1] = vc_o_4_4[2];
    data_i_5_4[1] = data_o_4_4[2];
    valid_i_5_4[1] = valid_o_4_4[2];
    ready_i_5_4[1] = ready_o_4_4[2];
    vc_i_5_4[0] = vc_i[5][4];
    data_i_5_4[0] = data_i[5][4];
    valid_i_5_4[0] = valid_i[5][4];
    ready_i_5_4[0] = ready_i[5][4];
end


/*Router 5,5*/    
cast_router #(
    .routing_table                  (routing_table_5_5)
)router_5_5(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_5_5),
    .data_i                         (data_i_5_5),
    .valid_i                        (valid_i_5_5),
    .ready_o                        (ready_o_5_5),
    .vc_o                           (vc_o_5_5),
    .data_o                         (data_o_5_5),
    .valid_o                        (valid_o_5_5),
    .ready_i                        (ready_i_5_5)
);


always_comb begin
    vc_i_5_5[3] = vc_o_5_4[4];
    data_i_5_5[3] = data_o_5_4[4];
    valid_i_5_5[3] = valid_o_5_4[4];
    ready_i_5_5[3] = ready_o_5_4[4];
    vc_i_5_5[4] = vc_o_5_6[3];
    data_i_5_5[4] = data_o_5_6[3];
    valid_i_5_5[4] = valid_o_5_6[3];
    ready_i_5_5[4] = ready_o_5_6[3];
    vc_i_5_5[1] = vc_o_4_5[2];
    data_i_5_5[1] = data_o_4_5[2];
    valid_i_5_5[1] = valid_o_4_5[2];
    ready_i_5_5[1] = ready_o_4_5[2];
    vc_i_5_5[0] = vc_i[5][5];
    data_i_5_5[0] = data_i[5][5];
    valid_i_5_5[0] = valid_i[5][5];
    ready_i_5_5[0] = ready_i[5][5];
end


/*Router 5,6*/    
cast_router #(
    .routing_table                  (routing_table_5_6)
)router_5_6(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_5_6),
    .data_i                         (data_i_5_6),
    .valid_i                        (valid_i_5_6),
    .ready_o                        (ready_o_5_6),
    .vc_o                           (vc_o_5_6),
    .data_o                         (data_o_5_6),
    .valid_o                        (valid_o_5_6),
    .ready_i                        (ready_i_5_6)
);


always_comb begin
    vc_i_5_6[3] = vc_o_5_5[4];
    data_i_5_6[3] = data_o_5_5[4];
    valid_i_5_6[3] = valid_o_5_5[4];
    ready_i_5_6[3] = ready_o_5_5[4];
    vc_i_5_6[4] = vc_o_5_7[3];
    data_i_5_6[4] = data_o_5_7[3];
    valid_i_5_6[4] = valid_o_5_7[3];
    ready_i_5_6[4] = ready_o_5_7[3];
    vc_i_5_6[1] = vc_o_4_6[2];
    data_i_5_6[1] = data_o_4_6[2];
    valid_i_5_6[1] = valid_o_4_6[2];
    ready_i_5_6[1] = ready_o_4_6[2];
    vc_i_5_6[0] = vc_i[5][6];
    data_i_5_6[0] = data_i[5][6];
    valid_i_5_6[0] = valid_i[5][6];
    ready_i_5_6[0] = ready_i[5][6];
end


/*Router 5,7*/    
cast_router #(
    .routing_table                  (routing_table_5_7)
)router_5_7(
    .clk                            (clk),
    .rstn                           (rstn),
    .vc_i                           (vc_i_5_7),
    .data_i                         (data_i_5_7),
    .valid_i                        (valid_i_5_7),
    .ready_o                        (ready_o_5_7),
    .vc_o                           (vc_o_5_7),
    .data_o                         (data_o_5_7),
    .valid_o                        (valid_o_5_7),
    .ready_i                        (ready_i_5_7)
);


always_comb begin
    vc_i_5_7[3] = vc_o_5_6[4];
    data_i_5_7[3] = data_o_5_6[4];
    valid_i_5_7[3] = valid_o_5_6[4];
    ready_i_5_7[3] = ready_o_5_6[4];
    vc_i_5_7[1] = vc_o_4_7[2];
    data_i_5_7[1] = data_o_4_7[2];
    valid_i_5_7[1] = valid_o_4_7[2];
    ready_i_5_7[1] = ready_o_4_7[2];
    vc_i_5_7[0] = vc_i[5][7];
    data_i_5_7[0] = data_i[5][7];
    valid_i_5_7[0] = valid_i[5][7];
    ready_i_5_7[0] = ready_i[5][7];
end


endmodule
