
`include "params.svh"
`include "connection_config.svh"

module system(
    input       wire                            clk,
    input       wire                            rstn,

    // inject ports
    input       wire        [`DW-1:0]           data_i_inject,
    input       wire                            valid_i_inject,
    output      wire                            ready_o_inject,

    // eject ports
    output      wire        [`DW-1:0]           data_o_eject [`EPN],
    output      wire                            valid_o_eject [`EPN],
    input       wire                            ready_i_eject [`EPN]
);

logic       [`DW-1:0]           cast_gather_data_t2n [`NW] [`NH];
logic                           cast_gather_valid_t2n [`NW] [`NH];
logic                           cast_gather_ready_n2t [`NW] [`NH];

logic       [`DW-1:0]           cast_data_n2t [`NW] [`NH];
logic                           cast_valid_n2t [`NW] [`NH];
logic                           cast_ready_t2n [`NW] [`NH];

logic       [`DW-1:0]           gather_data_n2t [`NW] [`NH];
logic                           gather_valid_n2t [`NW] [`NH];
logic                           gather_ready_t2n [`NW] [`NH];   

logic       [`DW-1:0]           merge_data_n2t [`NW] [`NH];
logic                           merge_valid_n2t [`NW] [`NH];
logic                           merge_ready_t2n [`NW] [`NH];

logic       [`DW-1:0]           merge_data_t2n [`NW] [`NH];
logic                           merge_valid_t2n [`NW] [`NH];
logic                           merge_ready_n2t [`NW] [`NH];

network network(
    .clk                                        (clk),
    .rstn                                       (rstn),

    .cast_gather_data_i                         (cast_gather_data_t2n),
    .cast_gather_valid_i                        (cast_gather_valid_t2n),
    .cast_gather_ready_o                        (cast_gather_ready_n2t),

    .cast_data_o                                (cast_data_n2t),
    .cast_valid_o                               (cast_valid_n2t),
    .cast_ready_i                               (cast_ready_t2n),      

    .gather_data_o                              (gather_data_n2t),
    .gather_valid_o                             (gather_valid_n2t),
    .gather_ready_i                             (gather_ready_t2n),

    .merge_data_i                               (merge_data_t2n),
    .merge_valid_i                              (merge_valid_t2n),
    .merge_ready_o                              (merge_ready_n2t),

    .merge_data_o                               (merge_data_n2t),
    .merge_valid_o                              (merge_valid_n2t),
    .merge_ready_i                              (merge_ready_t2n)
);


assign cast_ready_t2n[0][0] = 0;

virtual_tile #(
    .cast_out                       (cast_out[0][0]),
    .merge_in                       (merge_in[0][0]),
    .merge_out                      (merge_out[0][0]),
    .gather_in                      (gather_in[0][0]),
    .gather_out                     (gather_out[0][0]),
    .x                              (0),
    .y                              (0)
)tile_0_0(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (data_i_inject),
    .cast_valid_i                   (valid_i_inject),
    .cast_ready_o                   (ready_o_inject),

    // merge in
    .merge_data_i                   (merge_data_n2t[0][0]),
    .merge_valid_i                  (merge_valid_n2t[0][0]),
    .merge_ready_o                  (merge_ready_t2n[0][0]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[0][0]),
    .gather_valid_i                 (gather_valid_n2t[0][0]),
    .gather_ready_o                 (gather_ready_t2n[0][0]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[0][0]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[0][0]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[0][0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[0][0]),
    .merge_valid_o                  (merge_valid_t2n[0][0]),
    .merge_ready_i                  (merge_ready_n2t[0][0])
);


virtual_tile #(
    .cast_out                       (cast_out[0][1]),
    .merge_in                       (merge_in[0][1]),
    .merge_out                      (merge_out[0][1]),
    .gather_in                      (gather_in[0][1]),
    .gather_out                     (gather_out[0][1]),
    .x                              (0),
    .y                              (1)
)tile_0_1(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[0][1]),
    .cast_valid_i                   (cast_valid_n2t[0][1]),
    .cast_ready_o                   (cast_ready_t2n[0][1]),

    // merge in
    .merge_data_i                   (merge_data_n2t[0][1]),
    .merge_valid_i                  (merge_valid_n2t[0][1]),
    .merge_ready_o                  (merge_ready_t2n[0][1]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[0][1]),
    .gather_valid_i                 (gather_valid_n2t[0][1]),
    .gather_ready_o                 (gather_ready_t2n[0][1]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[0][1]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[0][1]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[0][1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[0][1]),
    .merge_valid_o                  (merge_valid_t2n[0][1]),
    .merge_ready_i                  (merge_ready_n2t[0][1])
);


virtual_tile #(
    .cast_out                       (cast_out[0][2]),
    .merge_in                       (merge_in[0][2]),
    .merge_out                      (merge_out[0][2]),
    .gather_in                      (gather_in[0][2]),
    .gather_out                     (gather_out[0][2]),
    .x                              (0),
    .y                              (2)
)tile_0_2(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[0][2]),
    .cast_valid_i                   (cast_valid_n2t[0][2]),
    .cast_ready_o                   (cast_ready_t2n[0][2]),

    // merge in
    .merge_data_i                   (merge_data_n2t[0][2]),
    .merge_valid_i                  (merge_valid_n2t[0][2]),
    .merge_ready_o                  (merge_ready_t2n[0][2]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[0][2]),
    .gather_valid_i                 (gather_valid_n2t[0][2]),
    .gather_ready_o                 (gather_ready_t2n[0][2]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[0][2]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[0][2]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[0][2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[0][2]),
    .merge_valid_o                  (merge_valid_t2n[0][2]),
    .merge_ready_i                  (merge_ready_n2t[0][2])
);


virtual_tile #(
    .cast_out                       (cast_out[0][3]),
    .merge_in                       (merge_in[0][3]),
    .merge_out                      (merge_out[0][3]),
    .gather_in                      (gather_in[0][3]),
    .gather_out                     (gather_out[0][3]),
    .x                              (0),
    .y                              (3)
)tile_0_3(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[0][3]),
    .cast_valid_i                   (cast_valid_n2t[0][3]),
    .cast_ready_o                   (cast_ready_t2n[0][3]),

    // merge in
    .merge_data_i                   (merge_data_n2t[0][3]),
    .merge_valid_i                  (merge_valid_n2t[0][3]),
    .merge_ready_o                  (merge_ready_t2n[0][3]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[0][3]),
    .gather_valid_i                 (gather_valid_n2t[0][3]),
    .gather_ready_o                 (gather_ready_t2n[0][3]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[0][3]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[0][3]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[0][3]),

    // merge out
    .merge_data_o                   (merge_data_t2n[0][3]),
    .merge_valid_o                  (merge_valid_t2n[0][3]),
    .merge_ready_i                  (merge_ready_n2t[0][3])
);


virtual_tile #(
    .cast_out                       (cast_out[0][4]),
    .merge_in                       (merge_in[0][4]),
    .merge_out                      (merge_out[0][4]),
    .gather_in                      (gather_in[0][4]),
    .gather_out                     (gather_out[0][4]),
    .x                              (0),
    .y                              (4)
)tile_0_4(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[0][4]),
    .cast_valid_i                   (cast_valid_n2t[0][4]),
    .cast_ready_o                   (cast_ready_t2n[0][4]),

    // merge in
    .merge_data_i                   (merge_data_n2t[0][4]),
    .merge_valid_i                  (merge_valid_n2t[0][4]),
    .merge_ready_o                  (merge_ready_t2n[0][4]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[0][4]),
    .gather_valid_i                 (gather_valid_n2t[0][4]),
    .gather_ready_o                 (gather_ready_t2n[0][4]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[0][4]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[0][4]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[0][4]),

    // merge out
    .merge_data_o                   (merge_data_t2n[0][4]),
    .merge_valid_o                  (merge_valid_t2n[0][4]),
    .merge_ready_i                  (merge_ready_n2t[0][4])
);


virtual_tile #(
    .cast_out                       (cast_out[0][5]),
    .merge_in                       (merge_in[0][5]),
    .merge_out                      (merge_out[0][5]),
    .gather_in                      (gather_in[0][5]),
    .gather_out                     (gather_out[0][5]),
    .x                              (0),
    .y                              (5)
)tile_0_5(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[0][5]),
    .cast_valid_i                   (cast_valid_n2t[0][5]),
    .cast_ready_o                   (cast_ready_t2n[0][5]),

    // merge in
    .merge_data_i                   (merge_data_n2t[0][5]),
    .merge_valid_i                  (merge_valid_n2t[0][5]),
    .merge_ready_o                  (merge_ready_t2n[0][5]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[0][5]),
    .gather_valid_i                 (gather_valid_n2t[0][5]),
    .gather_ready_o                 (gather_ready_t2n[0][5]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[0][5]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[0][5]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[0][5]),

    // merge out
    .merge_data_o                   (merge_data_t2n[0][5]),
    .merge_valid_o                  (merge_valid_t2n[0][5]),
    .merge_ready_i                  (merge_ready_n2t[0][5])
);


virtual_tile #(
    .cast_out                       (cast_out[0][6]),
    .merge_in                       (merge_in[0][6]),
    .merge_out                      (merge_out[0][6]),
    .gather_in                      (gather_in[0][6]),
    .gather_out                     (gather_out[0][6]),
    .x                              (0),
    .y                              (6)
)tile_0_6(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[0][6]),
    .cast_valid_i                   (cast_valid_n2t[0][6]),
    .cast_ready_o                   (cast_ready_t2n[0][6]),

    // merge in
    .merge_data_i                   (merge_data_n2t[0][6]),
    .merge_valid_i                  (merge_valid_n2t[0][6]),
    .merge_ready_o                  (merge_ready_t2n[0][6]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[0][6]),
    .gather_valid_i                 (gather_valid_n2t[0][6]),
    .gather_ready_o                 (gather_ready_t2n[0][6]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[0][6]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[0][6]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[0][6]),

    // merge out
    .merge_data_o                   (merge_data_t2n[0][6]),
    .merge_valid_o                  (merge_valid_t2n[0][6]),
    .merge_ready_i                  (merge_ready_n2t[0][6])
);


virtual_tile #(
    .cast_out                       (cast_out[0][7]),
    .merge_in                       (merge_in[0][7]),
    .merge_out                      (merge_out[0][7]),
    .gather_in                      (gather_in[0][7]),
    .gather_out                     (gather_out[0][7]),
    .x                              (0),
    .y                              (7)
)tile_0_7(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[0][7]),
    .cast_valid_i                   (cast_valid_n2t[0][7]),
    .cast_ready_o                   (cast_ready_t2n[0][7]),

    // merge in
    .merge_data_i                   (merge_data_n2t[0][7]),
    .merge_valid_i                  (merge_valid_n2t[0][7]),
    .merge_ready_o                  (merge_ready_t2n[0][7]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[0][7]),
    .gather_valid_i                 (gather_valid_n2t[0][7]),
    .gather_ready_o                 (gather_ready_t2n[0][7]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[0][7]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[0][7]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[0][7]),

    // merge out
    .merge_data_o                   (merge_data_t2n[0][7]),
    .merge_valid_o                  (merge_valid_t2n[0][7]),
    .merge_ready_i                  (merge_ready_n2t[0][7])
);


virtual_tile #(
    .cast_out                       (cast_out[0][8]),
    .merge_in                       (merge_in[0][8]),
    .merge_out                      (merge_out[0][8]),
    .gather_in                      (gather_in[0][8]),
    .gather_out                     (gather_out[0][8]),
    .x                              (0),
    .y                              (8)
)tile_0_8(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[0][8]),
    .cast_valid_i                   (cast_valid_n2t[0][8]),
    .cast_ready_o                   (cast_ready_t2n[0][8]),

    // merge in
    .merge_data_i                   (merge_data_n2t[0][8]),
    .merge_valid_i                  (merge_valid_n2t[0][8]),
    .merge_ready_o                  (merge_ready_t2n[0][8]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[0][8]),
    .gather_valid_i                 (gather_valid_n2t[0][8]),
    .gather_ready_o                 (gather_ready_t2n[0][8]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[0][8]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[0][8]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[0][8]),

    // merge out
    .merge_data_o                   (merge_data_t2n[0][8]),
    .merge_valid_o                  (merge_valid_t2n[0][8]),
    .merge_ready_i                  (merge_ready_n2t[0][8])
);


virtual_tile #(
    .cast_out                       (cast_out[1][0]),
    .merge_in                       (merge_in[1][0]),
    .merge_out                      (merge_out[1][0]),
    .gather_in                      (gather_in[1][0]),
    .gather_out                     (gather_out[1][0]),
    .x                              (1),
    .y                              (0)
)tile_1_0(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[1][0]),
    .cast_valid_i                   (cast_valid_n2t[1][0]),
    .cast_ready_o                   (cast_ready_t2n[1][0]),

    // merge in
    .merge_data_i                   (merge_data_n2t[1][0]),
    .merge_valid_i                  (merge_valid_n2t[1][0]),
    .merge_ready_o                  (merge_ready_t2n[1][0]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[1][0]),
    .gather_valid_i                 (gather_valid_n2t[1][0]),
    .gather_ready_o                 (gather_ready_t2n[1][0]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[1][0]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[1][0]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[1][0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[1][0]),
    .merge_valid_o                  (merge_valid_t2n[1][0]),
    .merge_ready_i                  (merge_ready_n2t[1][0])
);


virtual_tile #(
    .cast_out                       (cast_out[1][1]),
    .merge_in                       (merge_in[1][1]),
    .merge_out                      (merge_out[1][1]),
    .gather_in                      (gather_in[1][1]),
    .gather_out                     (gather_out[1][1]),
    .x                              (1),
    .y                              (1)
)tile_1_1(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[1][1]),
    .cast_valid_i                   (cast_valid_n2t[1][1]),
    .cast_ready_o                   (cast_ready_t2n[1][1]),

    // merge in
    .merge_data_i                   (merge_data_n2t[1][1]),
    .merge_valid_i                  (merge_valid_n2t[1][1]),
    .merge_ready_o                  (merge_ready_t2n[1][1]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[1][1]),
    .gather_valid_i                 (gather_valid_n2t[1][1]),
    .gather_ready_o                 (gather_ready_t2n[1][1]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[1][1]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[1][1]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[1][1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[1][1]),
    .merge_valid_o                  (merge_valid_t2n[1][1]),
    .merge_ready_i                  (merge_ready_n2t[1][1])
);


virtual_tile #(
    .cast_out                       (cast_out[1][2]),
    .merge_in                       (merge_in[1][2]),
    .merge_out                      (merge_out[1][2]),
    .gather_in                      (gather_in[1][2]),
    .gather_out                     (gather_out[1][2]),
    .x                              (1),
    .y                              (2)
)tile_1_2(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[1][2]),
    .cast_valid_i                   (cast_valid_n2t[1][2]),
    .cast_ready_o                   (cast_ready_t2n[1][2]),

    // merge in
    .merge_data_i                   (merge_data_n2t[1][2]),
    .merge_valid_i                  (merge_valid_n2t[1][2]),
    .merge_ready_o                  (merge_ready_t2n[1][2]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[1][2]),
    .gather_valid_i                 (gather_valid_n2t[1][2]),
    .gather_ready_o                 (gather_ready_t2n[1][2]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[1][2]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[1][2]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[1][2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[1][2]),
    .merge_valid_o                  (merge_valid_t2n[1][2]),
    .merge_ready_i                  (merge_ready_n2t[1][2])
);


virtual_tile #(
    .cast_out                       (cast_out[1][3]),
    .merge_in                       (merge_in[1][3]),
    .merge_out                      (merge_out[1][3]),
    .gather_in                      (gather_in[1][3]),
    .gather_out                     (gather_out[1][3]),
    .x                              (1),
    .y                              (3)
)tile_1_3(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[1][3]),
    .cast_valid_i                   (cast_valid_n2t[1][3]),
    .cast_ready_o                   (cast_ready_t2n[1][3]),

    // merge in
    .merge_data_i                   (merge_data_n2t[1][3]),
    .merge_valid_i                  (merge_valid_n2t[1][3]),
    .merge_ready_o                  (merge_ready_t2n[1][3]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[1][3]),
    .gather_valid_i                 (gather_valid_n2t[1][3]),
    .gather_ready_o                 (gather_ready_t2n[1][3]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[1][3]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[1][3]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[1][3]),

    // merge out
    .merge_data_o                   (merge_data_t2n[1][3]),
    .merge_valid_o                  (merge_valid_t2n[1][3]),
    .merge_ready_i                  (merge_ready_n2t[1][3])
);


virtual_tile #(
    .cast_out                       (cast_out[1][4]),
    .merge_in                       (merge_in[1][4]),
    .merge_out                      (merge_out[1][4]),
    .gather_in                      (gather_in[1][4]),
    .gather_out                     (gather_out[1][4]),
    .x                              (1),
    .y                              (4)
)tile_1_4(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[1][4]),
    .cast_valid_i                   (cast_valid_n2t[1][4]),
    .cast_ready_o                   (cast_ready_t2n[1][4]),

    // merge in
    .merge_data_i                   (merge_data_n2t[1][4]),
    .merge_valid_i                  (merge_valid_n2t[1][4]),
    .merge_ready_o                  (merge_ready_t2n[1][4]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[1][4]),
    .gather_valid_i                 (gather_valid_n2t[1][4]),
    .gather_ready_o                 (gather_ready_t2n[1][4]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[1][4]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[1][4]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[1][4]),

    // merge out
    .merge_data_o                   (merge_data_t2n[1][4]),
    .merge_valid_o                  (merge_valid_t2n[1][4]),
    .merge_ready_i                  (merge_ready_n2t[1][4])
);


virtual_tile #(
    .cast_out                       (cast_out[1][5]),
    .merge_in                       (merge_in[1][5]),
    .merge_out                      (merge_out[1][5]),
    .gather_in                      (gather_in[1][5]),
    .gather_out                     (gather_out[1][5]),
    .x                              (1),
    .y                              (5)
)tile_1_5(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[1][5]),
    .cast_valid_i                   (cast_valid_n2t[1][5]),
    .cast_ready_o                   (cast_ready_t2n[1][5]),

    // merge in
    .merge_data_i                   (merge_data_n2t[1][5]),
    .merge_valid_i                  (merge_valid_n2t[1][5]),
    .merge_ready_o                  (merge_ready_t2n[1][5]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[1][5]),
    .gather_valid_i                 (gather_valid_n2t[1][5]),
    .gather_ready_o                 (gather_ready_t2n[1][5]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[1][5]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[1][5]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[1][5]),

    // merge out
    .merge_data_o                   (merge_data_t2n[1][5]),
    .merge_valid_o                  (merge_valid_t2n[1][5]),
    .merge_ready_i                  (merge_ready_n2t[1][5])
);


virtual_tile #(
    .cast_out                       (cast_out[1][6]),
    .merge_in                       (merge_in[1][6]),
    .merge_out                      (merge_out[1][6]),
    .gather_in                      (gather_in[1][6]),
    .gather_out                     (gather_out[1][6]),
    .x                              (1),
    .y                              (6)
)tile_1_6(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[1][6]),
    .cast_valid_i                   (cast_valid_n2t[1][6]),
    .cast_ready_o                   (cast_ready_t2n[1][6]),

    // merge in
    .merge_data_i                   (merge_data_n2t[1][6]),
    .merge_valid_i                  (merge_valid_n2t[1][6]),
    .merge_ready_o                  (merge_ready_t2n[1][6]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[1][6]),
    .gather_valid_i                 (gather_valid_n2t[1][6]),
    .gather_ready_o                 (gather_ready_t2n[1][6]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[1][6]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[1][6]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[1][6]),

    // merge out
    .merge_data_o                   (merge_data_t2n[1][6]),
    .merge_valid_o                  (merge_valid_t2n[1][6]),
    .merge_ready_i                  (merge_ready_n2t[1][6])
);


virtual_tile #(
    .cast_out                       (cast_out[1][7]),
    .merge_in                       (merge_in[1][7]),
    .merge_out                      (merge_out[1][7]),
    .gather_in                      (gather_in[1][7]),
    .gather_out                     (gather_out[1][7]),
    .x                              (1),
    .y                              (7)
)tile_1_7(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[1][7]),
    .cast_valid_i                   (cast_valid_n2t[1][7]),
    .cast_ready_o                   (cast_ready_t2n[1][7]),

    // merge in
    .merge_data_i                   (merge_data_n2t[1][7]),
    .merge_valid_i                  (merge_valid_n2t[1][7]),
    .merge_ready_o                  (merge_ready_t2n[1][7]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[1][7]),
    .gather_valid_i                 (gather_valid_n2t[1][7]),
    .gather_ready_o                 (gather_ready_t2n[1][7]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[1][7]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[1][7]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[1][7]),

    // merge out
    .merge_data_o                   (merge_data_t2n[1][7]),
    .merge_valid_o                  (merge_valid_t2n[1][7]),
    .merge_ready_i                  (merge_ready_n2t[1][7])
);


virtual_tile #(
    .cast_out                       (cast_out[1][8]),
    .merge_in                       (merge_in[1][8]),
    .merge_out                      (merge_out[1][8]),
    .gather_in                      (gather_in[1][8]),
    .gather_out                     (gather_out[1][8]),
    .x                              (1),
    .y                              (8)
)tile_1_8(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[1][8]),
    .cast_valid_i                   (cast_valid_n2t[1][8]),
    .cast_ready_o                   (cast_ready_t2n[1][8]),

    // merge in
    .merge_data_i                   (merge_data_n2t[1][8]),
    .merge_valid_i                  (merge_valid_n2t[1][8]),
    .merge_ready_o                  (merge_ready_t2n[1][8]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[1][8]),
    .gather_valid_i                 (gather_valid_n2t[1][8]),
    .gather_ready_o                 (gather_ready_t2n[1][8]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[1][8]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[1][8]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[1][8]),

    // merge out
    .merge_data_o                   (merge_data_t2n[1][8]),
    .merge_valid_o                  (merge_valid_t2n[1][8]),
    .merge_ready_i                  (merge_ready_n2t[1][8])
);


virtual_tile #(
    .cast_out                       (cast_out[2][0]),
    .merge_in                       (merge_in[2][0]),
    .merge_out                      (merge_out[2][0]),
    .gather_in                      (gather_in[2][0]),
    .gather_out                     (gather_out[2][0]),
    .x                              (2),
    .y                              (0)
)tile_2_0(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[2][0]),
    .cast_valid_i                   (cast_valid_n2t[2][0]),
    .cast_ready_o                   (cast_ready_t2n[2][0]),

    // merge in
    .merge_data_i                   (merge_data_n2t[2][0]),
    .merge_valid_i                  (merge_valid_n2t[2][0]),
    .merge_ready_o                  (merge_ready_t2n[2][0]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[2][0]),
    .gather_valid_i                 (gather_valid_n2t[2][0]),
    .gather_ready_o                 (gather_ready_t2n[2][0]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[2][0]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[2][0]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[2][0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[2][0]),
    .merge_valid_o                  (merge_valid_t2n[2][0]),
    .merge_ready_i                  (merge_ready_n2t[2][0])
);


virtual_tile #(
    .cast_out                       (cast_out[2][1]),
    .merge_in                       (merge_in[2][1]),
    .merge_out                      (merge_out[2][1]),
    .gather_in                      (gather_in[2][1]),
    .gather_out                     (gather_out[2][1]),
    .x                              (2),
    .y                              (1)
)tile_2_1(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[2][1]),
    .cast_valid_i                   (cast_valid_n2t[2][1]),
    .cast_ready_o                   (cast_ready_t2n[2][1]),

    // merge in
    .merge_data_i                   (merge_data_n2t[2][1]),
    .merge_valid_i                  (merge_valid_n2t[2][1]),
    .merge_ready_o                  (merge_ready_t2n[2][1]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[2][1]),
    .gather_valid_i                 (gather_valid_n2t[2][1]),
    .gather_ready_o                 (gather_ready_t2n[2][1]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[2][1]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[2][1]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[2][1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[2][1]),
    .merge_valid_o                  (merge_valid_t2n[2][1]),
    .merge_ready_i                  (merge_ready_n2t[2][1])
);


virtual_tile #(
    .cast_out                       (cast_out[2][2]),
    .merge_in                       (merge_in[2][2]),
    .merge_out                      (merge_out[2][2]),
    .gather_in                      (gather_in[2][2]),
    .gather_out                     (gather_out[2][2]),
    .x                              (2),
    .y                              (2)
)tile_2_2(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[2][2]),
    .cast_valid_i                   (cast_valid_n2t[2][2]),
    .cast_ready_o                   (cast_ready_t2n[2][2]),

    // merge in
    .merge_data_i                   (merge_data_n2t[2][2]),
    .merge_valid_i                  (merge_valid_n2t[2][2]),
    .merge_ready_o                  (merge_ready_t2n[2][2]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[2][2]),
    .gather_valid_i                 (gather_valid_n2t[2][2]),
    .gather_ready_o                 (gather_ready_t2n[2][2]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[2][2]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[2][2]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[2][2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[2][2]),
    .merge_valid_o                  (merge_valid_t2n[2][2]),
    .merge_ready_i                  (merge_ready_n2t[2][2])
);


virtual_tile #(
    .cast_out                       (cast_out[2][3]),
    .merge_in                       (merge_in[2][3]),
    .merge_out                      (merge_out[2][3]),
    .gather_in                      (gather_in[2][3]),
    .gather_out                     (gather_out[2][3]),
    .x                              (2),
    .y                              (3)
)tile_2_3(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[2][3]),
    .cast_valid_i                   (cast_valid_n2t[2][3]),
    .cast_ready_o                   (cast_ready_t2n[2][3]),

    // merge in
    .merge_data_i                   (merge_data_n2t[2][3]),
    .merge_valid_i                  (merge_valid_n2t[2][3]),
    .merge_ready_o                  (merge_ready_t2n[2][3]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[2][3]),
    .gather_valid_i                 (gather_valid_n2t[2][3]),
    .gather_ready_o                 (gather_ready_t2n[2][3]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[2][3]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[2][3]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[2][3]),

    // merge out
    .merge_data_o                   (merge_data_t2n[2][3]),
    .merge_valid_o                  (merge_valid_t2n[2][3]),
    .merge_ready_i                  (merge_ready_n2t[2][3])
);


virtual_tile #(
    .cast_out                       (cast_out[2][4]),
    .merge_in                       (merge_in[2][4]),
    .merge_out                      (merge_out[2][4]),
    .gather_in                      (gather_in[2][4]),
    .gather_out                     (gather_out[2][4]),
    .x                              (2),
    .y                              (4)
)tile_2_4(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[2][4]),
    .cast_valid_i                   (cast_valid_n2t[2][4]),
    .cast_ready_o                   (cast_ready_t2n[2][4]),

    // merge in
    .merge_data_i                   (merge_data_n2t[2][4]),
    .merge_valid_i                  (merge_valid_n2t[2][4]),
    .merge_ready_o                  (merge_ready_t2n[2][4]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[2][4]),
    .gather_valid_i                 (gather_valid_n2t[2][4]),
    .gather_ready_o                 (gather_ready_t2n[2][4]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[2][4]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[2][4]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[2][4]),

    // merge out
    .merge_data_o                   (merge_data_t2n[2][4]),
    .merge_valid_o                  (merge_valid_t2n[2][4]),
    .merge_ready_i                  (merge_ready_n2t[2][4])
);


virtual_tile #(
    .cast_out                       (cast_out[2][5]),
    .merge_in                       (merge_in[2][5]),
    .merge_out                      (merge_out[2][5]),
    .gather_in                      (gather_in[2][5]),
    .gather_out                     (gather_out[2][5]),
    .x                              (2),
    .y                              (5)
)tile_2_5(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[2][5]),
    .cast_valid_i                   (cast_valid_n2t[2][5]),
    .cast_ready_o                   (cast_ready_t2n[2][5]),

    // merge in
    .merge_data_i                   (merge_data_n2t[2][5]),
    .merge_valid_i                  (merge_valid_n2t[2][5]),
    .merge_ready_o                  (merge_ready_t2n[2][5]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[2][5]),
    .gather_valid_i                 (gather_valid_n2t[2][5]),
    .gather_ready_o                 (gather_ready_t2n[2][5]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[2][5]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[2][5]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[2][5]),

    // merge out
    .merge_data_o                   (merge_data_t2n[2][5]),
    .merge_valid_o                  (merge_valid_t2n[2][5]),
    .merge_ready_i                  (merge_ready_n2t[2][5])
);


virtual_tile #(
    .cast_out                       (cast_out[2][6]),
    .merge_in                       (merge_in[2][6]),
    .merge_out                      (merge_out[2][6]),
    .gather_in                      (gather_in[2][6]),
    .gather_out                     (gather_out[2][6]),
    .x                              (2),
    .y                              (6)
)tile_2_6(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[2][6]),
    .cast_valid_i                   (cast_valid_n2t[2][6]),
    .cast_ready_o                   (cast_ready_t2n[2][6]),

    // merge in
    .merge_data_i                   (merge_data_n2t[2][6]),
    .merge_valid_i                  (merge_valid_n2t[2][6]),
    .merge_ready_o                  (merge_ready_t2n[2][6]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[2][6]),
    .gather_valid_i                 (gather_valid_n2t[2][6]),
    .gather_ready_o                 (gather_ready_t2n[2][6]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[2][6]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[2][6]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[2][6]),

    // merge out
    .merge_data_o                   (merge_data_t2n[2][6]),
    .merge_valid_o                  (merge_valid_t2n[2][6]),
    .merge_ready_i                  (merge_ready_n2t[2][6])
);


virtual_tile #(
    .cast_out                       (cast_out[2][7]),
    .merge_in                       (merge_in[2][7]),
    .merge_out                      (merge_out[2][7]),
    .gather_in                      (gather_in[2][7]),
    .gather_out                     (gather_out[2][7]),
    .x                              (2),
    .y                              (7)
)tile_2_7(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[2][7]),
    .cast_valid_i                   (cast_valid_n2t[2][7]),
    .cast_ready_o                   (cast_ready_t2n[2][7]),

    // merge in
    .merge_data_i                   (merge_data_n2t[2][7]),
    .merge_valid_i                  (merge_valid_n2t[2][7]),
    .merge_ready_o                  (merge_ready_t2n[2][7]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[2][7]),
    .gather_valid_i                 (gather_valid_n2t[2][7]),
    .gather_ready_o                 (gather_ready_t2n[2][7]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[2][7]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[2][7]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[2][7]),

    // merge out
    .merge_data_o                   (merge_data_t2n[2][7]),
    .merge_valid_o                  (merge_valid_t2n[2][7]),
    .merge_ready_i                  (merge_ready_n2t[2][7])
);


assign cast_gather_data_t2n[2][8] = 0;
assign cast_gather_valid_t2n[2][8] = 0;

virtual_tile #(
    .cast_out                       (cast_out[2][8]),
    .merge_in                       (merge_in[2][8]),
    .merge_out                      (merge_out[2][8]),
    .gather_in                      (gather_in[2][8]),
    .gather_out                     (gather_out[2][8]),
    .x                              (2),
    .y                              (8)
)tile_2_8(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[2][8]),
    .cast_valid_i                   (cast_valid_n2t[2][8]),
    .cast_ready_o                   (cast_ready_t2n[2][8]),

    // merge in
    .merge_data_i                   (merge_data_n2t[2][8]),
    .merge_valid_i                  (merge_valid_n2t[2][8]),
    .merge_ready_o                  (merge_ready_t2n[2][8]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[2][8]),
    .gather_valid_i                 (gather_valid_n2t[2][8]),
    .gather_ready_o                 (gather_ready_t2n[2][8]),

    // cast gather out
    .cast_gather_data_o             (data_o_eject[1]),
    .cast_gather_valid_o            (valid_o_eject[1]),   
    .cast_gather_ready_i            (ready_i_eject[1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[2][8]),
    .merge_valid_o                  (merge_valid_t2n[2][8]),
    .merge_ready_i                  (merge_ready_n2t[2][8])
);


virtual_tile #(
    .cast_out                       (cast_out[3][0]),
    .merge_in                       (merge_in[3][0]),
    .merge_out                      (merge_out[3][0]),
    .gather_in                      (gather_in[3][0]),
    .gather_out                     (gather_out[3][0]),
    .x                              (3),
    .y                              (0)
)tile_3_0(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[3][0]),
    .cast_valid_i                   (cast_valid_n2t[3][0]),
    .cast_ready_o                   (cast_ready_t2n[3][0]),

    // merge in
    .merge_data_i                   (merge_data_n2t[3][0]),
    .merge_valid_i                  (merge_valid_n2t[3][0]),
    .merge_ready_o                  (merge_ready_t2n[3][0]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[3][0]),
    .gather_valid_i                 (gather_valid_n2t[3][0]),
    .gather_ready_o                 (gather_ready_t2n[3][0]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[3][0]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[3][0]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[3][0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[3][0]),
    .merge_valid_o                  (merge_valid_t2n[3][0]),
    .merge_ready_i                  (merge_ready_n2t[3][0])
);


virtual_tile #(
    .cast_out                       (cast_out[3][1]),
    .merge_in                       (merge_in[3][1]),
    .merge_out                      (merge_out[3][1]),
    .gather_in                      (gather_in[3][1]),
    .gather_out                     (gather_out[3][1]),
    .x                              (3),
    .y                              (1)
)tile_3_1(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[3][1]),
    .cast_valid_i                   (cast_valid_n2t[3][1]),
    .cast_ready_o                   (cast_ready_t2n[3][1]),

    // merge in
    .merge_data_i                   (merge_data_n2t[3][1]),
    .merge_valid_i                  (merge_valid_n2t[3][1]),
    .merge_ready_o                  (merge_ready_t2n[3][1]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[3][1]),
    .gather_valid_i                 (gather_valid_n2t[3][1]),
    .gather_ready_o                 (gather_ready_t2n[3][1]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[3][1]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[3][1]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[3][1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[3][1]),
    .merge_valid_o                  (merge_valid_t2n[3][1]),
    .merge_ready_i                  (merge_ready_n2t[3][1])
);


virtual_tile #(
    .cast_out                       (cast_out[3][2]),
    .merge_in                       (merge_in[3][2]),
    .merge_out                      (merge_out[3][2]),
    .gather_in                      (gather_in[3][2]),
    .gather_out                     (gather_out[3][2]),
    .x                              (3),
    .y                              (2)
)tile_3_2(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[3][2]),
    .cast_valid_i                   (cast_valid_n2t[3][2]),
    .cast_ready_o                   (cast_ready_t2n[3][2]),

    // merge in
    .merge_data_i                   (merge_data_n2t[3][2]),
    .merge_valid_i                  (merge_valid_n2t[3][2]),
    .merge_ready_o                  (merge_ready_t2n[3][2]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[3][2]),
    .gather_valid_i                 (gather_valid_n2t[3][2]),
    .gather_ready_o                 (gather_ready_t2n[3][2]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[3][2]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[3][2]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[3][2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[3][2]),
    .merge_valid_o                  (merge_valid_t2n[3][2]),
    .merge_ready_i                  (merge_ready_n2t[3][2])
);


virtual_tile #(
    .cast_out                       (cast_out[3][3]),
    .merge_in                       (merge_in[3][3]),
    .merge_out                      (merge_out[3][3]),
    .gather_in                      (gather_in[3][3]),
    .gather_out                     (gather_out[3][3]),
    .x                              (3),
    .y                              (3)
)tile_3_3(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[3][3]),
    .cast_valid_i                   (cast_valid_n2t[3][3]),
    .cast_ready_o                   (cast_ready_t2n[3][3]),

    // merge in
    .merge_data_i                   (merge_data_n2t[3][3]),
    .merge_valid_i                  (merge_valid_n2t[3][3]),
    .merge_ready_o                  (merge_ready_t2n[3][3]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[3][3]),
    .gather_valid_i                 (gather_valid_n2t[3][3]),
    .gather_ready_o                 (gather_ready_t2n[3][3]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[3][3]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[3][3]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[3][3]),

    // merge out
    .merge_data_o                   (merge_data_t2n[3][3]),
    .merge_valid_o                  (merge_valid_t2n[3][3]),
    .merge_ready_i                  (merge_ready_n2t[3][3])
);


virtual_tile #(
    .cast_out                       (cast_out[3][4]),
    .merge_in                       (merge_in[3][4]),
    .merge_out                      (merge_out[3][4]),
    .gather_in                      (gather_in[3][4]),
    .gather_out                     (gather_out[3][4]),
    .x                              (3),
    .y                              (4)
)tile_3_4(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[3][4]),
    .cast_valid_i                   (cast_valid_n2t[3][4]),
    .cast_ready_o                   (cast_ready_t2n[3][4]),

    // merge in
    .merge_data_i                   (merge_data_n2t[3][4]),
    .merge_valid_i                  (merge_valid_n2t[3][4]),
    .merge_ready_o                  (merge_ready_t2n[3][4]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[3][4]),
    .gather_valid_i                 (gather_valid_n2t[3][4]),
    .gather_ready_o                 (gather_ready_t2n[3][4]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[3][4]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[3][4]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[3][4]),

    // merge out
    .merge_data_o                   (merge_data_t2n[3][4]),
    .merge_valid_o                  (merge_valid_t2n[3][4]),
    .merge_ready_i                  (merge_ready_n2t[3][4])
);


virtual_tile #(
    .cast_out                       (cast_out[3][5]),
    .merge_in                       (merge_in[3][5]),
    .merge_out                      (merge_out[3][5]),
    .gather_in                      (gather_in[3][5]),
    .gather_out                     (gather_out[3][5]),
    .x                              (3),
    .y                              (5)
)tile_3_5(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[3][5]),
    .cast_valid_i                   (cast_valid_n2t[3][5]),
    .cast_ready_o                   (cast_ready_t2n[3][5]),

    // merge in
    .merge_data_i                   (merge_data_n2t[3][5]),
    .merge_valid_i                  (merge_valid_n2t[3][5]),
    .merge_ready_o                  (merge_ready_t2n[3][5]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[3][5]),
    .gather_valid_i                 (gather_valid_n2t[3][5]),
    .gather_ready_o                 (gather_ready_t2n[3][5]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[3][5]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[3][5]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[3][5]),

    // merge out
    .merge_data_o                   (merge_data_t2n[3][5]),
    .merge_valid_o                  (merge_valid_t2n[3][5]),
    .merge_ready_i                  (merge_ready_n2t[3][5])
);


assign cast_gather_data_t2n[3][6] = 0;
assign cast_gather_valid_t2n[3][6] = 0;

virtual_tile #(
    .cast_out                       (cast_out[3][6]),
    .merge_in                       (merge_in[3][6]),
    .merge_out                      (merge_out[3][6]),
    .gather_in                      (gather_in[3][6]),
    .gather_out                     (gather_out[3][6]),
    .x                              (3),
    .y                              (6)
)tile_3_6(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[3][6]),
    .cast_valid_i                   (cast_valid_n2t[3][6]),
    .cast_ready_o                   (cast_ready_t2n[3][6]),

    // merge in
    .merge_data_i                   (merge_data_n2t[3][6]),
    .merge_valid_i                  (merge_valid_n2t[3][6]),
    .merge_ready_o                  (merge_ready_t2n[3][6]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[3][6]),
    .gather_valid_i                 (gather_valid_n2t[3][6]),
    .gather_ready_o                 (gather_ready_t2n[3][6]),

    // cast gather out
    .cast_gather_data_o             (data_o_eject[0]),
    .cast_gather_valid_o            (valid_o_eject[0]),   
    .cast_gather_ready_i            (ready_i_eject[0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[3][6]),
    .merge_valid_o                  (merge_valid_t2n[3][6]),
    .merge_ready_i                  (merge_ready_n2t[3][6])
);


virtual_tile #(
    .cast_out                       (cast_out[3][7]),
    .merge_in                       (merge_in[3][7]),
    .merge_out                      (merge_out[3][7]),
    .gather_in                      (gather_in[3][7]),
    .gather_out                     (gather_out[3][7]),
    .x                              (3),
    .y                              (7)
)tile_3_7(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[3][7]),
    .cast_valid_i                   (cast_valid_n2t[3][7]),
    .cast_ready_o                   (cast_ready_t2n[3][7]),

    // merge in
    .merge_data_i                   (merge_data_n2t[3][7]),
    .merge_valid_i                  (merge_valid_n2t[3][7]),
    .merge_ready_o                  (merge_ready_t2n[3][7]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[3][7]),
    .gather_valid_i                 (gather_valid_n2t[3][7]),
    .gather_ready_o                 (gather_ready_t2n[3][7]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[3][7]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[3][7]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[3][7]),

    // merge out
    .merge_data_o                   (merge_data_t2n[3][7]),
    .merge_valid_o                  (merge_valid_t2n[3][7]),
    .merge_ready_i                  (merge_ready_n2t[3][7])
);


virtual_tile #(
    .cast_out                       (cast_out[3][8]),
    .merge_in                       (merge_in[3][8]),
    .merge_out                      (merge_out[3][8]),
    .gather_in                      (gather_in[3][8]),
    .gather_out                     (gather_out[3][8]),
    .x                              (3),
    .y                              (8)
)tile_3_8(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[3][8]),
    .cast_valid_i                   (cast_valid_n2t[3][8]),
    .cast_ready_o                   (cast_ready_t2n[3][8]),

    // merge in
    .merge_data_i                   (merge_data_n2t[3][8]),
    .merge_valid_i                  (merge_valid_n2t[3][8]),
    .merge_ready_o                  (merge_ready_t2n[3][8]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[3][8]),
    .gather_valid_i                 (gather_valid_n2t[3][8]),
    .gather_ready_o                 (gather_ready_t2n[3][8]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[3][8]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[3][8]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[3][8]),

    // merge out
    .merge_data_o                   (merge_data_t2n[3][8]),
    .merge_valid_o                  (merge_valid_t2n[3][8]),
    .merge_ready_i                  (merge_ready_n2t[3][8])
);


virtual_tile #(
    .cast_out                       (cast_out[4][0]),
    .merge_in                       (merge_in[4][0]),
    .merge_out                      (merge_out[4][0]),
    .gather_in                      (gather_in[4][0]),
    .gather_out                     (gather_out[4][0]),
    .x                              (4),
    .y                              (0)
)tile_4_0(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[4][0]),
    .cast_valid_i                   (cast_valid_n2t[4][0]),
    .cast_ready_o                   (cast_ready_t2n[4][0]),

    // merge in
    .merge_data_i                   (merge_data_n2t[4][0]),
    .merge_valid_i                  (merge_valid_n2t[4][0]),
    .merge_ready_o                  (merge_ready_t2n[4][0]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[4][0]),
    .gather_valid_i                 (gather_valid_n2t[4][0]),
    .gather_ready_o                 (gather_ready_t2n[4][0]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[4][0]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[4][0]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[4][0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[4][0]),
    .merge_valid_o                  (merge_valid_t2n[4][0]),
    .merge_ready_i                  (merge_ready_n2t[4][0])
);


virtual_tile #(
    .cast_out                       (cast_out[4][1]),
    .merge_in                       (merge_in[4][1]),
    .merge_out                      (merge_out[4][1]),
    .gather_in                      (gather_in[4][1]),
    .gather_out                     (gather_out[4][1]),
    .x                              (4),
    .y                              (1)
)tile_4_1(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[4][1]),
    .cast_valid_i                   (cast_valid_n2t[4][1]),
    .cast_ready_o                   (cast_ready_t2n[4][1]),

    // merge in
    .merge_data_i                   (merge_data_n2t[4][1]),
    .merge_valid_i                  (merge_valid_n2t[4][1]),
    .merge_ready_o                  (merge_ready_t2n[4][1]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[4][1]),
    .gather_valid_i                 (gather_valid_n2t[4][1]),
    .gather_ready_o                 (gather_ready_t2n[4][1]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[4][1]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[4][1]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[4][1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[4][1]),
    .merge_valid_o                  (merge_valid_t2n[4][1]),
    .merge_ready_i                  (merge_ready_n2t[4][1])
);


virtual_tile #(
    .cast_out                       (cast_out[4][2]),
    .merge_in                       (merge_in[4][2]),
    .merge_out                      (merge_out[4][2]),
    .gather_in                      (gather_in[4][2]),
    .gather_out                     (gather_out[4][2]),
    .x                              (4),
    .y                              (2)
)tile_4_2(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[4][2]),
    .cast_valid_i                   (cast_valid_n2t[4][2]),
    .cast_ready_o                   (cast_ready_t2n[4][2]),

    // merge in
    .merge_data_i                   (merge_data_n2t[4][2]),
    .merge_valid_i                  (merge_valid_n2t[4][2]),
    .merge_ready_o                  (merge_ready_t2n[4][2]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[4][2]),
    .gather_valid_i                 (gather_valid_n2t[4][2]),
    .gather_ready_o                 (gather_ready_t2n[4][2]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[4][2]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[4][2]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[4][2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[4][2]),
    .merge_valid_o                  (merge_valid_t2n[4][2]),
    .merge_ready_i                  (merge_ready_n2t[4][2])
);


virtual_tile #(
    .cast_out                       (cast_out[4][3]),
    .merge_in                       (merge_in[4][3]),
    .merge_out                      (merge_out[4][3]),
    .gather_in                      (gather_in[4][3]),
    .gather_out                     (gather_out[4][3]),
    .x                              (4),
    .y                              (3)
)tile_4_3(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[4][3]),
    .cast_valid_i                   (cast_valid_n2t[4][3]),
    .cast_ready_o                   (cast_ready_t2n[4][3]),

    // merge in
    .merge_data_i                   (merge_data_n2t[4][3]),
    .merge_valid_i                  (merge_valid_n2t[4][3]),
    .merge_ready_o                  (merge_ready_t2n[4][3]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[4][3]),
    .gather_valid_i                 (gather_valid_n2t[4][3]),
    .gather_ready_o                 (gather_ready_t2n[4][3]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[4][3]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[4][3]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[4][3]),

    // merge out
    .merge_data_o                   (merge_data_t2n[4][3]),
    .merge_valid_o                  (merge_valid_t2n[4][3]),
    .merge_ready_i                  (merge_ready_n2t[4][3])
);


virtual_tile #(
    .cast_out                       (cast_out[4][4]),
    .merge_in                       (merge_in[4][4]),
    .merge_out                      (merge_out[4][4]),
    .gather_in                      (gather_in[4][4]),
    .gather_out                     (gather_out[4][4]),
    .x                              (4),
    .y                              (4)
)tile_4_4(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[4][4]),
    .cast_valid_i                   (cast_valid_n2t[4][4]),
    .cast_ready_o                   (cast_ready_t2n[4][4]),

    // merge in
    .merge_data_i                   (merge_data_n2t[4][4]),
    .merge_valid_i                  (merge_valid_n2t[4][4]),
    .merge_ready_o                  (merge_ready_t2n[4][4]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[4][4]),
    .gather_valid_i                 (gather_valid_n2t[4][4]),
    .gather_ready_o                 (gather_ready_t2n[4][4]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[4][4]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[4][4]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[4][4]),

    // merge out
    .merge_data_o                   (merge_data_t2n[4][4]),
    .merge_valid_o                  (merge_valid_t2n[4][4]),
    .merge_ready_i                  (merge_ready_n2t[4][4])
);


virtual_tile #(
    .cast_out                       (cast_out[4][5]),
    .merge_in                       (merge_in[4][5]),
    .merge_out                      (merge_out[4][5]),
    .gather_in                      (gather_in[4][5]),
    .gather_out                     (gather_out[4][5]),
    .x                              (4),
    .y                              (5)
)tile_4_5(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[4][5]),
    .cast_valid_i                   (cast_valid_n2t[4][5]),
    .cast_ready_o                   (cast_ready_t2n[4][5]),

    // merge in
    .merge_data_i                   (merge_data_n2t[4][5]),
    .merge_valid_i                  (merge_valid_n2t[4][5]),
    .merge_ready_o                  (merge_ready_t2n[4][5]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[4][5]),
    .gather_valid_i                 (gather_valid_n2t[4][5]),
    .gather_ready_o                 (gather_ready_t2n[4][5]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[4][5]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[4][5]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[4][5]),

    // merge out
    .merge_data_o                   (merge_data_t2n[4][5]),
    .merge_valid_o                  (merge_valid_t2n[4][5]),
    .merge_ready_i                  (merge_ready_n2t[4][5])
);


virtual_tile #(
    .cast_out                       (cast_out[4][6]),
    .merge_in                       (merge_in[4][6]),
    .merge_out                      (merge_out[4][6]),
    .gather_in                      (gather_in[4][6]),
    .gather_out                     (gather_out[4][6]),
    .x                              (4),
    .y                              (6)
)tile_4_6(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[4][6]),
    .cast_valid_i                   (cast_valid_n2t[4][6]),
    .cast_ready_o                   (cast_ready_t2n[4][6]),

    // merge in
    .merge_data_i                   (merge_data_n2t[4][6]),
    .merge_valid_i                  (merge_valid_n2t[4][6]),
    .merge_ready_o                  (merge_ready_t2n[4][6]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[4][6]),
    .gather_valid_i                 (gather_valid_n2t[4][6]),
    .gather_ready_o                 (gather_ready_t2n[4][6]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[4][6]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[4][6]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[4][6]),

    // merge out
    .merge_data_o                   (merge_data_t2n[4][6]),
    .merge_valid_o                  (merge_valid_t2n[4][6]),
    .merge_ready_i                  (merge_ready_n2t[4][6])
);


virtual_tile #(
    .cast_out                       (cast_out[4][7]),
    .merge_in                       (merge_in[4][7]),
    .merge_out                      (merge_out[4][7]),
    .gather_in                      (gather_in[4][7]),
    .gather_out                     (gather_out[4][7]),
    .x                              (4),
    .y                              (7)
)tile_4_7(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[4][7]),
    .cast_valid_i                   (cast_valid_n2t[4][7]),
    .cast_ready_o                   (cast_ready_t2n[4][7]),

    // merge in
    .merge_data_i                   (merge_data_n2t[4][7]),
    .merge_valid_i                  (merge_valid_n2t[4][7]),
    .merge_ready_o                  (merge_ready_t2n[4][7]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[4][7]),
    .gather_valid_i                 (gather_valid_n2t[4][7]),
    .gather_ready_o                 (gather_ready_t2n[4][7]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[4][7]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[4][7]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[4][7]),

    // merge out
    .merge_data_o                   (merge_data_t2n[4][7]),
    .merge_valid_o                  (merge_valid_t2n[4][7]),
    .merge_ready_i                  (merge_ready_n2t[4][7])
);


virtual_tile #(
    .cast_out                       (cast_out[4][8]),
    .merge_in                       (merge_in[4][8]),
    .merge_out                      (merge_out[4][8]),
    .gather_in                      (gather_in[4][8]),
    .gather_out                     (gather_out[4][8]),
    .x                              (4),
    .y                              (8)
)tile_4_8(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[4][8]),
    .cast_valid_i                   (cast_valid_n2t[4][8]),
    .cast_ready_o                   (cast_ready_t2n[4][8]),

    // merge in
    .merge_data_i                   (merge_data_n2t[4][8]),
    .merge_valid_i                  (merge_valid_n2t[4][8]),
    .merge_ready_o                  (merge_ready_t2n[4][8]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[4][8]),
    .gather_valid_i                 (gather_valid_n2t[4][8]),
    .gather_ready_o                 (gather_ready_t2n[4][8]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[4][8]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[4][8]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[4][8]),

    // merge out
    .merge_data_o                   (merge_data_t2n[4][8]),
    .merge_valid_o                  (merge_valid_t2n[4][8]),
    .merge_ready_i                  (merge_ready_n2t[4][8])
);


virtual_tile #(
    .cast_out                       (cast_out[5][0]),
    .merge_in                       (merge_in[5][0]),
    .merge_out                      (merge_out[5][0]),
    .gather_in                      (gather_in[5][0]),
    .gather_out                     (gather_out[5][0]),
    .x                              (5),
    .y                              (0)
)tile_5_0(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[5][0]),
    .cast_valid_i                   (cast_valid_n2t[5][0]),
    .cast_ready_o                   (cast_ready_t2n[5][0]),

    // merge in
    .merge_data_i                   (merge_data_n2t[5][0]),
    .merge_valid_i                  (merge_valid_n2t[5][0]),
    .merge_ready_o                  (merge_ready_t2n[5][0]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[5][0]),
    .gather_valid_i                 (gather_valid_n2t[5][0]),
    .gather_ready_o                 (gather_ready_t2n[5][0]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[5][0]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[5][0]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[5][0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[5][0]),
    .merge_valid_o                  (merge_valid_t2n[5][0]),
    .merge_ready_i                  (merge_ready_n2t[5][0])
);


virtual_tile #(
    .cast_out                       (cast_out[5][1]),
    .merge_in                       (merge_in[5][1]),
    .merge_out                      (merge_out[5][1]),
    .gather_in                      (gather_in[5][1]),
    .gather_out                     (gather_out[5][1]),
    .x                              (5),
    .y                              (1)
)tile_5_1(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[5][1]),
    .cast_valid_i                   (cast_valid_n2t[5][1]),
    .cast_ready_o                   (cast_ready_t2n[5][1]),

    // merge in
    .merge_data_i                   (merge_data_n2t[5][1]),
    .merge_valid_i                  (merge_valid_n2t[5][1]),
    .merge_ready_o                  (merge_ready_t2n[5][1]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[5][1]),
    .gather_valid_i                 (gather_valid_n2t[5][1]),
    .gather_ready_o                 (gather_ready_t2n[5][1]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[5][1]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[5][1]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[5][1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[5][1]),
    .merge_valid_o                  (merge_valid_t2n[5][1]),
    .merge_ready_i                  (merge_ready_n2t[5][1])
);


virtual_tile #(
    .cast_out                       (cast_out[5][2]),
    .merge_in                       (merge_in[5][2]),
    .merge_out                      (merge_out[5][2]),
    .gather_in                      (gather_in[5][2]),
    .gather_out                     (gather_out[5][2]),
    .x                              (5),
    .y                              (2)
)tile_5_2(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[5][2]),
    .cast_valid_i                   (cast_valid_n2t[5][2]),
    .cast_ready_o                   (cast_ready_t2n[5][2]),

    // merge in
    .merge_data_i                   (merge_data_n2t[5][2]),
    .merge_valid_i                  (merge_valid_n2t[5][2]),
    .merge_ready_o                  (merge_ready_t2n[5][2]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[5][2]),
    .gather_valid_i                 (gather_valid_n2t[5][2]),
    .gather_ready_o                 (gather_ready_t2n[5][2]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[5][2]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[5][2]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[5][2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[5][2]),
    .merge_valid_o                  (merge_valid_t2n[5][2]),
    .merge_ready_i                  (merge_ready_n2t[5][2])
);


virtual_tile #(
    .cast_out                       (cast_out[5][3]),
    .merge_in                       (merge_in[5][3]),
    .merge_out                      (merge_out[5][3]),
    .gather_in                      (gather_in[5][3]),
    .gather_out                     (gather_out[5][3]),
    .x                              (5),
    .y                              (3)
)tile_5_3(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[5][3]),
    .cast_valid_i                   (cast_valid_n2t[5][3]),
    .cast_ready_o                   (cast_ready_t2n[5][3]),

    // merge in
    .merge_data_i                   (merge_data_n2t[5][3]),
    .merge_valid_i                  (merge_valid_n2t[5][3]),
    .merge_ready_o                  (merge_ready_t2n[5][3]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[5][3]),
    .gather_valid_i                 (gather_valid_n2t[5][3]),
    .gather_ready_o                 (gather_ready_t2n[5][3]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[5][3]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[5][3]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[5][3]),

    // merge out
    .merge_data_o                   (merge_data_t2n[5][3]),
    .merge_valid_o                  (merge_valid_t2n[5][3]),
    .merge_ready_i                  (merge_ready_n2t[5][3])
);


virtual_tile #(
    .cast_out                       (cast_out[5][4]),
    .merge_in                       (merge_in[5][4]),
    .merge_out                      (merge_out[5][4]),
    .gather_in                      (gather_in[5][4]),
    .gather_out                     (gather_out[5][4]),
    .x                              (5),
    .y                              (4)
)tile_5_4(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[5][4]),
    .cast_valid_i                   (cast_valid_n2t[5][4]),
    .cast_ready_o                   (cast_ready_t2n[5][4]),

    // merge in
    .merge_data_i                   (merge_data_n2t[5][4]),
    .merge_valid_i                  (merge_valid_n2t[5][4]),
    .merge_ready_o                  (merge_ready_t2n[5][4]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[5][4]),
    .gather_valid_i                 (gather_valid_n2t[5][4]),
    .gather_ready_o                 (gather_ready_t2n[5][4]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[5][4]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[5][4]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[5][4]),

    // merge out
    .merge_data_o                   (merge_data_t2n[5][4]),
    .merge_valid_o                  (merge_valid_t2n[5][4]),
    .merge_ready_i                  (merge_ready_n2t[5][4])
);


virtual_tile #(
    .cast_out                       (cast_out[5][5]),
    .merge_in                       (merge_in[5][5]),
    .merge_out                      (merge_out[5][5]),
    .gather_in                      (gather_in[5][5]),
    .gather_out                     (gather_out[5][5]),
    .x                              (5),
    .y                              (5)
)tile_5_5(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[5][5]),
    .cast_valid_i                   (cast_valid_n2t[5][5]),
    .cast_ready_o                   (cast_ready_t2n[5][5]),

    // merge in
    .merge_data_i                   (merge_data_n2t[5][5]),
    .merge_valid_i                  (merge_valid_n2t[5][5]),
    .merge_ready_o                  (merge_ready_t2n[5][5]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[5][5]),
    .gather_valid_i                 (gather_valid_n2t[5][5]),
    .gather_ready_o                 (gather_ready_t2n[5][5]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[5][5]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[5][5]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[5][5]),

    // merge out
    .merge_data_o                   (merge_data_t2n[5][5]),
    .merge_valid_o                  (merge_valid_t2n[5][5]),
    .merge_ready_i                  (merge_ready_n2t[5][5])
);


virtual_tile #(
    .cast_out                       (cast_out[5][6]),
    .merge_in                       (merge_in[5][6]),
    .merge_out                      (merge_out[5][6]),
    .gather_in                      (gather_in[5][6]),
    .gather_out                     (gather_out[5][6]),
    .x                              (5),
    .y                              (6)
)tile_5_6(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[5][6]),
    .cast_valid_i                   (cast_valid_n2t[5][6]),
    .cast_ready_o                   (cast_ready_t2n[5][6]),

    // merge in
    .merge_data_i                   (merge_data_n2t[5][6]),
    .merge_valid_i                  (merge_valid_n2t[5][6]),
    .merge_ready_o                  (merge_ready_t2n[5][6]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[5][6]),
    .gather_valid_i                 (gather_valid_n2t[5][6]),
    .gather_ready_o                 (gather_ready_t2n[5][6]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[5][6]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[5][6]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[5][6]),

    // merge out
    .merge_data_o                   (merge_data_t2n[5][6]),
    .merge_valid_o                  (merge_valid_t2n[5][6]),
    .merge_ready_i                  (merge_ready_n2t[5][6])
);


virtual_tile #(
    .cast_out                       (cast_out[5][7]),
    .merge_in                       (merge_in[5][7]),
    .merge_out                      (merge_out[5][7]),
    .gather_in                      (gather_in[5][7]),
    .gather_out                     (gather_out[5][7]),
    .x                              (5),
    .y                              (7)
)tile_5_7(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[5][7]),
    .cast_valid_i                   (cast_valid_n2t[5][7]),
    .cast_ready_o                   (cast_ready_t2n[5][7]),

    // merge in
    .merge_data_i                   (merge_data_n2t[5][7]),
    .merge_valid_i                  (merge_valid_n2t[5][7]),
    .merge_ready_o                  (merge_ready_t2n[5][7]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[5][7]),
    .gather_valid_i                 (gather_valid_n2t[5][7]),
    .gather_ready_o                 (gather_ready_t2n[5][7]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[5][7]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[5][7]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[5][7]),

    // merge out
    .merge_data_o                   (merge_data_t2n[5][7]),
    .merge_valid_o                  (merge_valid_t2n[5][7]),
    .merge_ready_i                  (merge_ready_n2t[5][7])
);


assign cast_gather_data_t2n[5][8] = 0;
assign cast_gather_valid_t2n[5][8] = 0;

virtual_tile #(
    .cast_out                       (cast_out[5][8]),
    .merge_in                       (merge_in[5][8]),
    .merge_out                      (merge_out[5][8]),
    .gather_in                      (gather_in[5][8]),
    .gather_out                     (gather_out[5][8]),
    .x                              (5),
    .y                              (8)
)tile_5_8(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[5][8]),
    .cast_valid_i                   (cast_valid_n2t[5][8]),
    .cast_ready_o                   (cast_ready_t2n[5][8]),

    // merge in
    .merge_data_i                   (merge_data_n2t[5][8]),
    .merge_valid_i                  (merge_valid_n2t[5][8]),
    .merge_ready_o                  (merge_ready_t2n[5][8]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[5][8]),
    .gather_valid_i                 (gather_valid_n2t[5][8]),
    .gather_ready_o                 (gather_ready_t2n[5][8]),

    // cast gather out
    .cast_gather_data_o             (data_o_eject[2]),
    .cast_gather_valid_o            (valid_o_eject[2]),   
    .cast_gather_ready_i            (ready_i_eject[2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[5][8]),
    .merge_valid_o                  (merge_valid_t2n[5][8]),
    .merge_ready_i                  (merge_ready_n2t[5][8])
);


virtual_tile #(
    .cast_out                       (cast_out[6][0]),
    .merge_in                       (merge_in[6][0]),
    .merge_out                      (merge_out[6][0]),
    .gather_in                      (gather_in[6][0]),
    .gather_out                     (gather_out[6][0]),
    .x                              (6),
    .y                              (0)
)tile_6_0(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[6][0]),
    .cast_valid_i                   (cast_valid_n2t[6][0]),
    .cast_ready_o                   (cast_ready_t2n[6][0]),

    // merge in
    .merge_data_i                   (merge_data_n2t[6][0]),
    .merge_valid_i                  (merge_valid_n2t[6][0]),
    .merge_ready_o                  (merge_ready_t2n[6][0]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[6][0]),
    .gather_valid_i                 (gather_valid_n2t[6][0]),
    .gather_ready_o                 (gather_ready_t2n[6][0]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[6][0]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[6][0]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[6][0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[6][0]),
    .merge_valid_o                  (merge_valid_t2n[6][0]),
    .merge_ready_i                  (merge_ready_n2t[6][0])
);


virtual_tile #(
    .cast_out                       (cast_out[6][1]),
    .merge_in                       (merge_in[6][1]),
    .merge_out                      (merge_out[6][1]),
    .gather_in                      (gather_in[6][1]),
    .gather_out                     (gather_out[6][1]),
    .x                              (6),
    .y                              (1)
)tile_6_1(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[6][1]),
    .cast_valid_i                   (cast_valid_n2t[6][1]),
    .cast_ready_o                   (cast_ready_t2n[6][1]),

    // merge in
    .merge_data_i                   (merge_data_n2t[6][1]),
    .merge_valid_i                  (merge_valid_n2t[6][1]),
    .merge_ready_o                  (merge_ready_t2n[6][1]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[6][1]),
    .gather_valid_i                 (gather_valid_n2t[6][1]),
    .gather_ready_o                 (gather_ready_t2n[6][1]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[6][1]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[6][1]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[6][1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[6][1]),
    .merge_valid_o                  (merge_valid_t2n[6][1]),
    .merge_ready_i                  (merge_ready_n2t[6][1])
);


virtual_tile #(
    .cast_out                       (cast_out[6][2]),
    .merge_in                       (merge_in[6][2]),
    .merge_out                      (merge_out[6][2]),
    .gather_in                      (gather_in[6][2]),
    .gather_out                     (gather_out[6][2]),
    .x                              (6),
    .y                              (2)
)tile_6_2(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[6][2]),
    .cast_valid_i                   (cast_valid_n2t[6][2]),
    .cast_ready_o                   (cast_ready_t2n[6][2]),

    // merge in
    .merge_data_i                   (merge_data_n2t[6][2]),
    .merge_valid_i                  (merge_valid_n2t[6][2]),
    .merge_ready_o                  (merge_ready_t2n[6][2]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[6][2]),
    .gather_valid_i                 (gather_valid_n2t[6][2]),
    .gather_ready_o                 (gather_ready_t2n[6][2]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[6][2]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[6][2]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[6][2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[6][2]),
    .merge_valid_o                  (merge_valid_t2n[6][2]),
    .merge_ready_i                  (merge_ready_n2t[6][2])
);


virtual_tile #(
    .cast_out                       (cast_out[6][3]),
    .merge_in                       (merge_in[6][3]),
    .merge_out                      (merge_out[6][3]),
    .gather_in                      (gather_in[6][3]),
    .gather_out                     (gather_out[6][3]),
    .x                              (6),
    .y                              (3)
)tile_6_3(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[6][3]),
    .cast_valid_i                   (cast_valid_n2t[6][3]),
    .cast_ready_o                   (cast_ready_t2n[6][3]),

    // merge in
    .merge_data_i                   (merge_data_n2t[6][3]),
    .merge_valid_i                  (merge_valid_n2t[6][3]),
    .merge_ready_o                  (merge_ready_t2n[6][3]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[6][3]),
    .gather_valid_i                 (gather_valid_n2t[6][3]),
    .gather_ready_o                 (gather_ready_t2n[6][3]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[6][3]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[6][3]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[6][3]),

    // merge out
    .merge_data_o                   (merge_data_t2n[6][3]),
    .merge_valid_o                  (merge_valid_t2n[6][3]),
    .merge_ready_i                  (merge_ready_n2t[6][3])
);


virtual_tile #(
    .cast_out                       (cast_out[6][4]),
    .merge_in                       (merge_in[6][4]),
    .merge_out                      (merge_out[6][4]),
    .gather_in                      (gather_in[6][4]),
    .gather_out                     (gather_out[6][4]),
    .x                              (6),
    .y                              (4)
)tile_6_4(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[6][4]),
    .cast_valid_i                   (cast_valid_n2t[6][4]),
    .cast_ready_o                   (cast_ready_t2n[6][4]),

    // merge in
    .merge_data_i                   (merge_data_n2t[6][4]),
    .merge_valid_i                  (merge_valid_n2t[6][4]),
    .merge_ready_o                  (merge_ready_t2n[6][4]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[6][4]),
    .gather_valid_i                 (gather_valid_n2t[6][4]),
    .gather_ready_o                 (gather_ready_t2n[6][4]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[6][4]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[6][4]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[6][4]),

    // merge out
    .merge_data_o                   (merge_data_t2n[6][4]),
    .merge_valid_o                  (merge_valid_t2n[6][4]),
    .merge_ready_i                  (merge_ready_n2t[6][4])
);


virtual_tile #(
    .cast_out                       (cast_out[6][5]),
    .merge_in                       (merge_in[6][5]),
    .merge_out                      (merge_out[6][5]),
    .gather_in                      (gather_in[6][5]),
    .gather_out                     (gather_out[6][5]),
    .x                              (6),
    .y                              (5)
)tile_6_5(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[6][5]),
    .cast_valid_i                   (cast_valid_n2t[6][5]),
    .cast_ready_o                   (cast_ready_t2n[6][5]),

    // merge in
    .merge_data_i                   (merge_data_n2t[6][5]),
    .merge_valid_i                  (merge_valid_n2t[6][5]),
    .merge_ready_o                  (merge_ready_t2n[6][5]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[6][5]),
    .gather_valid_i                 (gather_valid_n2t[6][5]),
    .gather_ready_o                 (gather_ready_t2n[6][5]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[6][5]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[6][5]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[6][5]),

    // merge out
    .merge_data_o                   (merge_data_t2n[6][5]),
    .merge_valid_o                  (merge_valid_t2n[6][5]),
    .merge_ready_i                  (merge_ready_n2t[6][5])
);


virtual_tile #(
    .cast_out                       (cast_out[6][6]),
    .merge_in                       (merge_in[6][6]),
    .merge_out                      (merge_out[6][6]),
    .gather_in                      (gather_in[6][6]),
    .gather_out                     (gather_out[6][6]),
    .x                              (6),
    .y                              (6)
)tile_6_6(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[6][6]),
    .cast_valid_i                   (cast_valid_n2t[6][6]),
    .cast_ready_o                   (cast_ready_t2n[6][6]),

    // merge in
    .merge_data_i                   (merge_data_n2t[6][6]),
    .merge_valid_i                  (merge_valid_n2t[6][6]),
    .merge_ready_o                  (merge_ready_t2n[6][6]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[6][6]),
    .gather_valid_i                 (gather_valid_n2t[6][6]),
    .gather_ready_o                 (gather_ready_t2n[6][6]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[6][6]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[6][6]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[6][6]),

    // merge out
    .merge_data_o                   (merge_data_t2n[6][6]),
    .merge_valid_o                  (merge_valid_t2n[6][6]),
    .merge_ready_i                  (merge_ready_n2t[6][6])
);


virtual_tile #(
    .cast_out                       (cast_out[6][7]),
    .merge_in                       (merge_in[6][7]),
    .merge_out                      (merge_out[6][7]),
    .gather_in                      (gather_in[6][7]),
    .gather_out                     (gather_out[6][7]),
    .x                              (6),
    .y                              (7)
)tile_6_7(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[6][7]),
    .cast_valid_i                   (cast_valid_n2t[6][7]),
    .cast_ready_o                   (cast_ready_t2n[6][7]),

    // merge in
    .merge_data_i                   (merge_data_n2t[6][7]),
    .merge_valid_i                  (merge_valid_n2t[6][7]),
    .merge_ready_o                  (merge_ready_t2n[6][7]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[6][7]),
    .gather_valid_i                 (gather_valid_n2t[6][7]),
    .gather_ready_o                 (gather_ready_t2n[6][7]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[6][7]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[6][7]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[6][7]),

    // merge out
    .merge_data_o                   (merge_data_t2n[6][7]),
    .merge_valid_o                  (merge_valid_t2n[6][7]),
    .merge_ready_i                  (merge_ready_n2t[6][7])
);


virtual_tile #(
    .cast_out                       (cast_out[6][8]),
    .merge_in                       (merge_in[6][8]),
    .merge_out                      (merge_out[6][8]),
    .gather_in                      (gather_in[6][8]),
    .gather_out                     (gather_out[6][8]),
    .x                              (6),
    .y                              (8)
)tile_6_8(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[6][8]),
    .cast_valid_i                   (cast_valid_n2t[6][8]),
    .cast_ready_o                   (cast_ready_t2n[6][8]),

    // merge in
    .merge_data_i                   (merge_data_n2t[6][8]),
    .merge_valid_i                  (merge_valid_n2t[6][8]),
    .merge_ready_o                  (merge_ready_t2n[6][8]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[6][8]),
    .gather_valid_i                 (gather_valid_n2t[6][8]),
    .gather_ready_o                 (gather_ready_t2n[6][8]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[6][8]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[6][8]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[6][8]),

    // merge out
    .merge_data_o                   (merge_data_t2n[6][8]),
    .merge_valid_o                  (merge_valid_t2n[6][8]),
    .merge_ready_i                  (merge_ready_n2t[6][8])
);


virtual_tile #(
    .cast_out                       (cast_out[7][0]),
    .merge_in                       (merge_in[7][0]),
    .merge_out                      (merge_out[7][0]),
    .gather_in                      (gather_in[7][0]),
    .gather_out                     (gather_out[7][0]),
    .x                              (7),
    .y                              (0)
)tile_7_0(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[7][0]),
    .cast_valid_i                   (cast_valid_n2t[7][0]),
    .cast_ready_o                   (cast_ready_t2n[7][0]),

    // merge in
    .merge_data_i                   (merge_data_n2t[7][0]),
    .merge_valid_i                  (merge_valid_n2t[7][0]),
    .merge_ready_o                  (merge_ready_t2n[7][0]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[7][0]),
    .gather_valid_i                 (gather_valid_n2t[7][0]),
    .gather_ready_o                 (gather_ready_t2n[7][0]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[7][0]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[7][0]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[7][0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[7][0]),
    .merge_valid_o                  (merge_valid_t2n[7][0]),
    .merge_ready_i                  (merge_ready_n2t[7][0])
);


virtual_tile #(
    .cast_out                       (cast_out[7][1]),
    .merge_in                       (merge_in[7][1]),
    .merge_out                      (merge_out[7][1]),
    .gather_in                      (gather_in[7][1]),
    .gather_out                     (gather_out[7][1]),
    .x                              (7),
    .y                              (1)
)tile_7_1(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[7][1]),
    .cast_valid_i                   (cast_valid_n2t[7][1]),
    .cast_ready_o                   (cast_ready_t2n[7][1]),

    // merge in
    .merge_data_i                   (merge_data_n2t[7][1]),
    .merge_valid_i                  (merge_valid_n2t[7][1]),
    .merge_ready_o                  (merge_ready_t2n[7][1]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[7][1]),
    .gather_valid_i                 (gather_valid_n2t[7][1]),
    .gather_ready_o                 (gather_ready_t2n[7][1]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[7][1]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[7][1]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[7][1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[7][1]),
    .merge_valid_o                  (merge_valid_t2n[7][1]),
    .merge_ready_i                  (merge_ready_n2t[7][1])
);


virtual_tile #(
    .cast_out                       (cast_out[7][2]),
    .merge_in                       (merge_in[7][2]),
    .merge_out                      (merge_out[7][2]),
    .gather_in                      (gather_in[7][2]),
    .gather_out                     (gather_out[7][2]),
    .x                              (7),
    .y                              (2)
)tile_7_2(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[7][2]),
    .cast_valid_i                   (cast_valid_n2t[7][2]),
    .cast_ready_o                   (cast_ready_t2n[7][2]),

    // merge in
    .merge_data_i                   (merge_data_n2t[7][2]),
    .merge_valid_i                  (merge_valid_n2t[7][2]),
    .merge_ready_o                  (merge_ready_t2n[7][2]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[7][2]),
    .gather_valid_i                 (gather_valid_n2t[7][2]),
    .gather_ready_o                 (gather_ready_t2n[7][2]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[7][2]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[7][2]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[7][2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[7][2]),
    .merge_valid_o                  (merge_valid_t2n[7][2]),
    .merge_ready_i                  (merge_ready_n2t[7][2])
);


virtual_tile #(
    .cast_out                       (cast_out[7][3]),
    .merge_in                       (merge_in[7][3]),
    .merge_out                      (merge_out[7][3]),
    .gather_in                      (gather_in[7][3]),
    .gather_out                     (gather_out[7][3]),
    .x                              (7),
    .y                              (3)
)tile_7_3(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[7][3]),
    .cast_valid_i                   (cast_valid_n2t[7][3]),
    .cast_ready_o                   (cast_ready_t2n[7][3]),

    // merge in
    .merge_data_i                   (merge_data_n2t[7][3]),
    .merge_valid_i                  (merge_valid_n2t[7][3]),
    .merge_ready_o                  (merge_ready_t2n[7][3]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[7][3]),
    .gather_valid_i                 (gather_valid_n2t[7][3]),
    .gather_ready_o                 (gather_ready_t2n[7][3]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[7][3]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[7][3]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[7][3]),

    // merge out
    .merge_data_o                   (merge_data_t2n[7][3]),
    .merge_valid_o                  (merge_valid_t2n[7][3]),
    .merge_ready_i                  (merge_ready_n2t[7][3])
);


virtual_tile #(
    .cast_out                       (cast_out[7][4]),
    .merge_in                       (merge_in[7][4]),
    .merge_out                      (merge_out[7][4]),
    .gather_in                      (gather_in[7][4]),
    .gather_out                     (gather_out[7][4]),
    .x                              (7),
    .y                              (4)
)tile_7_4(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[7][4]),
    .cast_valid_i                   (cast_valid_n2t[7][4]),
    .cast_ready_o                   (cast_ready_t2n[7][4]),

    // merge in
    .merge_data_i                   (merge_data_n2t[7][4]),
    .merge_valid_i                  (merge_valid_n2t[7][4]),
    .merge_ready_o                  (merge_ready_t2n[7][4]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[7][4]),
    .gather_valid_i                 (gather_valid_n2t[7][4]),
    .gather_ready_o                 (gather_ready_t2n[7][4]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[7][4]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[7][4]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[7][4]),

    // merge out
    .merge_data_o                   (merge_data_t2n[7][4]),
    .merge_valid_o                  (merge_valid_t2n[7][4]),
    .merge_ready_i                  (merge_ready_n2t[7][4])
);


virtual_tile #(
    .cast_out                       (cast_out[7][5]),
    .merge_in                       (merge_in[7][5]),
    .merge_out                      (merge_out[7][5]),
    .gather_in                      (gather_in[7][5]),
    .gather_out                     (gather_out[7][5]),
    .x                              (7),
    .y                              (5)
)tile_7_5(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[7][5]),
    .cast_valid_i                   (cast_valid_n2t[7][5]),
    .cast_ready_o                   (cast_ready_t2n[7][5]),

    // merge in
    .merge_data_i                   (merge_data_n2t[7][5]),
    .merge_valid_i                  (merge_valid_n2t[7][5]),
    .merge_ready_o                  (merge_ready_t2n[7][5]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[7][5]),
    .gather_valid_i                 (gather_valid_n2t[7][5]),
    .gather_ready_o                 (gather_ready_t2n[7][5]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[7][5]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[7][5]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[7][5]),

    // merge out
    .merge_data_o                   (merge_data_t2n[7][5]),
    .merge_valid_o                  (merge_valid_t2n[7][5]),
    .merge_ready_i                  (merge_ready_n2t[7][5])
);


virtual_tile #(
    .cast_out                       (cast_out[7][6]),
    .merge_in                       (merge_in[7][6]),
    .merge_out                      (merge_out[7][6]),
    .gather_in                      (gather_in[7][6]),
    .gather_out                     (gather_out[7][6]),
    .x                              (7),
    .y                              (6)
)tile_7_6(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[7][6]),
    .cast_valid_i                   (cast_valid_n2t[7][6]),
    .cast_ready_o                   (cast_ready_t2n[7][6]),

    // merge in
    .merge_data_i                   (merge_data_n2t[7][6]),
    .merge_valid_i                  (merge_valid_n2t[7][6]),
    .merge_ready_o                  (merge_ready_t2n[7][6]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[7][6]),
    .gather_valid_i                 (gather_valid_n2t[7][6]),
    .gather_ready_o                 (gather_ready_t2n[7][6]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[7][6]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[7][6]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[7][6]),

    // merge out
    .merge_data_o                   (merge_data_t2n[7][6]),
    .merge_valid_o                  (merge_valid_t2n[7][6]),
    .merge_ready_i                  (merge_ready_n2t[7][6])
);


virtual_tile #(
    .cast_out                       (cast_out[7][7]),
    .merge_in                       (merge_in[7][7]),
    .merge_out                      (merge_out[7][7]),
    .gather_in                      (gather_in[7][7]),
    .gather_out                     (gather_out[7][7]),
    .x                              (7),
    .y                              (7)
)tile_7_7(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[7][7]),
    .cast_valid_i                   (cast_valid_n2t[7][7]),
    .cast_ready_o                   (cast_ready_t2n[7][7]),

    // merge in
    .merge_data_i                   (merge_data_n2t[7][7]),
    .merge_valid_i                  (merge_valid_n2t[7][7]),
    .merge_ready_o                  (merge_ready_t2n[7][7]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[7][7]),
    .gather_valid_i                 (gather_valid_n2t[7][7]),
    .gather_ready_o                 (gather_ready_t2n[7][7]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[7][7]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[7][7]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[7][7]),

    // merge out
    .merge_data_o                   (merge_data_t2n[7][7]),
    .merge_valid_o                  (merge_valid_t2n[7][7]),
    .merge_ready_i                  (merge_ready_n2t[7][7])
);


virtual_tile #(
    .cast_out                       (cast_out[7][8]),
    .merge_in                       (merge_in[7][8]),
    .merge_out                      (merge_out[7][8]),
    .gather_in                      (gather_in[7][8]),
    .gather_out                     (gather_out[7][8]),
    .x                              (7),
    .y                              (8)
)tile_7_8(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[7][8]),
    .cast_valid_i                   (cast_valid_n2t[7][8]),
    .cast_ready_o                   (cast_ready_t2n[7][8]),

    // merge in
    .merge_data_i                   (merge_data_n2t[7][8]),
    .merge_valid_i                  (merge_valid_n2t[7][8]),
    .merge_ready_o                  (merge_ready_t2n[7][8]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[7][8]),
    .gather_valid_i                 (gather_valid_n2t[7][8]),
    .gather_ready_o                 (gather_ready_t2n[7][8]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[7][8]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[7][8]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[7][8]),

    // merge out
    .merge_data_o                   (merge_data_t2n[7][8]),
    .merge_valid_o                  (merge_valid_t2n[7][8]),
    .merge_ready_i                  (merge_ready_n2t[7][8])
);


virtual_tile #(
    .cast_out                       (cast_out[8][0]),
    .merge_in                       (merge_in[8][0]),
    .merge_out                      (merge_out[8][0]),
    .gather_in                      (gather_in[8][0]),
    .gather_out                     (gather_out[8][0]),
    .x                              (8),
    .y                              (0)
)tile_8_0(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[8][0]),
    .cast_valid_i                   (cast_valid_n2t[8][0]),
    .cast_ready_o                   (cast_ready_t2n[8][0]),

    // merge in
    .merge_data_i                   (merge_data_n2t[8][0]),
    .merge_valid_i                  (merge_valid_n2t[8][0]),
    .merge_ready_o                  (merge_ready_t2n[8][0]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[8][0]),
    .gather_valid_i                 (gather_valid_n2t[8][0]),
    .gather_ready_o                 (gather_ready_t2n[8][0]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[8][0]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[8][0]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[8][0]),

    // merge out
    .merge_data_o                   (merge_data_t2n[8][0]),
    .merge_valid_o                  (merge_valid_t2n[8][0]),
    .merge_ready_i                  (merge_ready_n2t[8][0])
);


virtual_tile #(
    .cast_out                       (cast_out[8][1]),
    .merge_in                       (merge_in[8][1]),
    .merge_out                      (merge_out[8][1]),
    .gather_in                      (gather_in[8][1]),
    .gather_out                     (gather_out[8][1]),
    .x                              (8),
    .y                              (1)
)tile_8_1(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[8][1]),
    .cast_valid_i                   (cast_valid_n2t[8][1]),
    .cast_ready_o                   (cast_ready_t2n[8][1]),

    // merge in
    .merge_data_i                   (merge_data_n2t[8][1]),
    .merge_valid_i                  (merge_valid_n2t[8][1]),
    .merge_ready_o                  (merge_ready_t2n[8][1]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[8][1]),
    .gather_valid_i                 (gather_valid_n2t[8][1]),
    .gather_ready_o                 (gather_ready_t2n[8][1]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[8][1]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[8][1]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[8][1]),

    // merge out
    .merge_data_o                   (merge_data_t2n[8][1]),
    .merge_valid_o                  (merge_valid_t2n[8][1]),
    .merge_ready_i                  (merge_ready_n2t[8][1])
);


virtual_tile #(
    .cast_out                       (cast_out[8][2]),
    .merge_in                       (merge_in[8][2]),
    .merge_out                      (merge_out[8][2]),
    .gather_in                      (gather_in[8][2]),
    .gather_out                     (gather_out[8][2]),
    .x                              (8),
    .y                              (2)
)tile_8_2(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[8][2]),
    .cast_valid_i                   (cast_valid_n2t[8][2]),
    .cast_ready_o                   (cast_ready_t2n[8][2]),

    // merge in
    .merge_data_i                   (merge_data_n2t[8][2]),
    .merge_valid_i                  (merge_valid_n2t[8][2]),
    .merge_ready_o                  (merge_ready_t2n[8][2]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[8][2]),
    .gather_valid_i                 (gather_valid_n2t[8][2]),
    .gather_ready_o                 (gather_ready_t2n[8][2]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[8][2]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[8][2]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[8][2]),

    // merge out
    .merge_data_o                   (merge_data_t2n[8][2]),
    .merge_valid_o                  (merge_valid_t2n[8][2]),
    .merge_ready_i                  (merge_ready_n2t[8][2])
);


virtual_tile #(
    .cast_out                       (cast_out[8][3]),
    .merge_in                       (merge_in[8][3]),
    .merge_out                      (merge_out[8][3]),
    .gather_in                      (gather_in[8][3]),
    .gather_out                     (gather_out[8][3]),
    .x                              (8),
    .y                              (3)
)tile_8_3(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[8][3]),
    .cast_valid_i                   (cast_valid_n2t[8][3]),
    .cast_ready_o                   (cast_ready_t2n[8][3]),

    // merge in
    .merge_data_i                   (merge_data_n2t[8][3]),
    .merge_valid_i                  (merge_valid_n2t[8][3]),
    .merge_ready_o                  (merge_ready_t2n[8][3]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[8][3]),
    .gather_valid_i                 (gather_valid_n2t[8][3]),
    .gather_ready_o                 (gather_ready_t2n[8][3]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[8][3]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[8][3]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[8][3]),

    // merge out
    .merge_data_o                   (merge_data_t2n[8][3]),
    .merge_valid_o                  (merge_valid_t2n[8][3]),
    .merge_ready_i                  (merge_ready_n2t[8][3])
);


virtual_tile #(
    .cast_out                       (cast_out[8][4]),
    .merge_in                       (merge_in[8][4]),
    .merge_out                      (merge_out[8][4]),
    .gather_in                      (gather_in[8][4]),
    .gather_out                     (gather_out[8][4]),
    .x                              (8),
    .y                              (4)
)tile_8_4(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[8][4]),
    .cast_valid_i                   (cast_valid_n2t[8][4]),
    .cast_ready_o                   (cast_ready_t2n[8][4]),

    // merge in
    .merge_data_i                   (merge_data_n2t[8][4]),
    .merge_valid_i                  (merge_valid_n2t[8][4]),
    .merge_ready_o                  (merge_ready_t2n[8][4]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[8][4]),
    .gather_valid_i                 (gather_valid_n2t[8][4]),
    .gather_ready_o                 (gather_ready_t2n[8][4]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[8][4]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[8][4]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[8][4]),

    // merge out
    .merge_data_o                   (merge_data_t2n[8][4]),
    .merge_valid_o                  (merge_valid_t2n[8][4]),
    .merge_ready_i                  (merge_ready_n2t[8][4])
);


virtual_tile #(
    .cast_out                       (cast_out[8][5]),
    .merge_in                       (merge_in[8][5]),
    .merge_out                      (merge_out[8][5]),
    .gather_in                      (gather_in[8][5]),
    .gather_out                     (gather_out[8][5]),
    .x                              (8),
    .y                              (5)
)tile_8_5(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[8][5]),
    .cast_valid_i                   (cast_valid_n2t[8][5]),
    .cast_ready_o                   (cast_ready_t2n[8][5]),

    // merge in
    .merge_data_i                   (merge_data_n2t[8][5]),
    .merge_valid_i                  (merge_valid_n2t[8][5]),
    .merge_ready_o                  (merge_ready_t2n[8][5]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[8][5]),
    .gather_valid_i                 (gather_valid_n2t[8][5]),
    .gather_ready_o                 (gather_ready_t2n[8][5]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[8][5]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[8][5]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[8][5]),

    // merge out
    .merge_data_o                   (merge_data_t2n[8][5]),
    .merge_valid_o                  (merge_valid_t2n[8][5]),
    .merge_ready_i                  (merge_ready_n2t[8][5])
);


virtual_tile #(
    .cast_out                       (cast_out[8][6]),
    .merge_in                       (merge_in[8][6]),
    .merge_out                      (merge_out[8][6]),
    .gather_in                      (gather_in[8][6]),
    .gather_out                     (gather_out[8][6]),
    .x                              (8),
    .y                              (6)
)tile_8_6(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[8][6]),
    .cast_valid_i                   (cast_valid_n2t[8][6]),
    .cast_ready_o                   (cast_ready_t2n[8][6]),

    // merge in
    .merge_data_i                   (merge_data_n2t[8][6]),
    .merge_valid_i                  (merge_valid_n2t[8][6]),
    .merge_ready_o                  (merge_ready_t2n[8][6]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[8][6]),
    .gather_valid_i                 (gather_valid_n2t[8][6]),
    .gather_ready_o                 (gather_ready_t2n[8][6]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[8][6]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[8][6]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[8][6]),

    // merge out
    .merge_data_o                   (merge_data_t2n[8][6]),
    .merge_valid_o                  (merge_valid_t2n[8][6]),
    .merge_ready_i                  (merge_ready_n2t[8][6])
);


virtual_tile #(
    .cast_out                       (cast_out[8][7]),
    .merge_in                       (merge_in[8][7]),
    .merge_out                      (merge_out[8][7]),
    .gather_in                      (gather_in[8][7]),
    .gather_out                     (gather_out[8][7]),
    .x                              (8),
    .y                              (7)
)tile_8_7(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[8][7]),
    .cast_valid_i                   (cast_valid_n2t[8][7]),
    .cast_ready_o                   (cast_ready_t2n[8][7]),

    // merge in
    .merge_data_i                   (merge_data_n2t[8][7]),
    .merge_valid_i                  (merge_valid_n2t[8][7]),
    .merge_ready_o                  (merge_ready_t2n[8][7]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[8][7]),
    .gather_valid_i                 (gather_valid_n2t[8][7]),
    .gather_ready_o                 (gather_ready_t2n[8][7]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[8][7]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[8][7]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[8][7]),

    // merge out
    .merge_data_o                   (merge_data_t2n[8][7]),
    .merge_valid_o                  (merge_valid_t2n[8][7]),
    .merge_ready_i                  (merge_ready_n2t[8][7])
);


virtual_tile #(
    .cast_out                       (cast_out[8][8]),
    .merge_in                       (merge_in[8][8]),
    .merge_out                      (merge_out[8][8]),
    .gather_in                      (gather_in[8][8]),
    .gather_out                     (gather_out[8][8]),
    .x                              (8),
    .y                              (8)
)tile_8_8(
    .clk                            (clk),
    .rstn                           (rstn), 

    // cast in
    .cast_data_i                    (cast_data_n2t[8][8]),
    .cast_valid_i                   (cast_valid_n2t[8][8]),
    .cast_ready_o                   (cast_ready_t2n[8][8]),

    // merge in
    .merge_data_i                   (merge_data_n2t[8][8]),
    .merge_valid_i                  (merge_valid_n2t[8][8]),
    .merge_ready_o                  (merge_ready_t2n[8][8]),

    // gather in 
    .gather_data_i                  (gather_data_n2t[8][8]),
    .gather_valid_i                 (gather_valid_n2t[8][8]),
    .gather_ready_o                 (gather_ready_t2n[8][8]),

    // cast gather out
    .cast_gather_data_o             (cast_gather_data_t2n[8][8]),
    .cast_gather_valid_o            (cast_gather_valid_t2n[8][8]),   
    .cast_gather_ready_i            (cast_gather_ready_n2t[8][8]),

    // merge out
    .merge_data_o                   (merge_data_t2n[8][8]),
    .merge_valid_o                  (merge_valid_t2n[8][8]),
    .merge_ready_i                  (merge_ready_n2t[8][8])
);


endmodule
